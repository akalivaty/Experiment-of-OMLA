

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793;

  OR2_X1 U372 ( .A1(n764), .A2(n490), .ZN(n491) );
  AND2_X1 U373 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U374 ( .A(n528), .B(n527), .ZN(n509) );
  XNOR2_X1 U375 ( .A(n355), .B(n354), .ZN(n771) );
  INV_X1 U376 ( .A(G128), .ZN(n507) );
  INV_X1 U377 ( .A(G104), .ZN(n356) );
  AND2_X2 U378 ( .A1(n720), .A2(n719), .ZN(n600) );
  XNOR2_X1 U379 ( .A(G143), .B(G104), .ZN(n553) );
  XNOR2_X1 U380 ( .A(G113), .B(KEYINPUT69), .ZN(n357) );
  OR2_X1 U381 ( .A1(n674), .A2(n414), .ZN(n359) );
  XNOR2_X1 U382 ( .A(G119), .B(G128), .ZN(n571) );
  XNOR2_X1 U383 ( .A(n405), .B(G472), .ZN(n725) );
  XOR2_X1 U384 ( .A(n502), .B(KEYINPUT41), .Z(n351) );
  XOR2_X1 U385 ( .A(KEYINPUT13), .B(G475), .Z(n352) );
  XNOR2_X2 U386 ( .A(n484), .B(n509), .ZN(n674) );
  NOR2_X2 U387 ( .A1(n723), .A2(n722), .ZN(n720) );
  NAND2_X2 U388 ( .A1(n360), .A2(n359), .ZN(n644) );
  AND2_X2 U389 ( .A1(n787), .A2(KEYINPUT44), .ZN(n468) );
  XNOR2_X2 U390 ( .A(n528), .B(n515), .ZN(n545) );
  INV_X4 U391 ( .A(G146), .ZN(n466) );
  INV_X1 U392 ( .A(KEYINPUT1), .ZN(n397) );
  NAND2_X1 U393 ( .A1(n377), .A2(n374), .ZN(n791) );
  NAND2_X1 U394 ( .A1(n376), .A2(n375), .ZN(n374) );
  AND2_X1 U395 ( .A1(n380), .A2(n378), .ZN(n377) );
  INV_X1 U396 ( .A(n733), .ZN(n376) );
  NAND2_X1 U397 ( .A1(n386), .A2(n383), .ZN(n733) );
  NOR2_X1 U398 ( .A1(n640), .A2(n389), .ZN(n375) );
  AND2_X1 U399 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U400 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U401 ( .A1(n398), .A2(n397), .ZN(n396) );
  OR2_X1 U402 ( .A1(n751), .A2(G902), .ZN(n372) );
  OR2_X1 U403 ( .A1(n669), .A2(G902), .ZN(n405) );
  OR2_X1 U404 ( .A1(n747), .A2(n399), .ZN(n398) );
  INV_X1 U405 ( .A(n414), .ZN(n366) );
  NAND2_X1 U406 ( .A1(G469), .A2(G902), .ZN(n403) );
  INV_X1 U407 ( .A(G469), .ZN(n401) );
  INV_X1 U408 ( .A(G119), .ZN(n392) );
  INV_X2 U409 ( .A(G953), .ZN(n781) );
  INV_X1 U410 ( .A(G902), .ZN(n400) );
  AND2_X1 U411 ( .A1(n492), .A2(n495), .ZN(n498) );
  INV_X1 U412 ( .A(n665), .ZN(n659) );
  OR2_X1 U413 ( .A1(n665), .A2(n664), .ZN(n666) );
  AND2_X1 U414 ( .A1(n634), .A2(n478), .ZN(n499) );
  XNOR2_X1 U415 ( .A(KEYINPUT32), .B(n591), .ZN(n788) );
  XNOR2_X1 U416 ( .A(n464), .B(n422), .ZN(n785) );
  XNOR2_X1 U417 ( .A(n453), .B(KEYINPUT31), .ZN(n456) );
  XNOR2_X1 U418 ( .A(n639), .B(n638), .ZN(n657) );
  XNOR2_X1 U419 ( .A(n426), .B(KEYINPUT96), .ZN(n599) );
  OR2_X1 U420 ( .A1(n711), .A2(n709), .ZN(n503) );
  XNOR2_X1 U421 ( .A(n616), .B(KEYINPUT28), .ZN(n617) );
  NAND2_X2 U422 ( .A1(n394), .A2(n393), .ZN(n719) );
  NOR2_X1 U423 ( .A1(n722), .A2(n615), .ZN(n643) );
  XNOR2_X1 U424 ( .A(n559), .B(KEYINPUT105), .ZN(n711) );
  NAND2_X1 U425 ( .A1(n395), .A2(KEYINPUT1), .ZN(n393) );
  NOR2_X1 U426 ( .A1(n603), .A2(n595), .ZN(n697) );
  AND2_X1 U427 ( .A1(n363), .A2(n361), .ZN(n360) );
  NAND2_X1 U428 ( .A1(n402), .A2(n398), .ZN(n395) );
  XNOR2_X1 U429 ( .A(n372), .B(n352), .ZN(n602) );
  XNOR2_X1 U430 ( .A(n485), .B(n486), .ZN(n484) );
  BUF_X1 U431 ( .A(n457), .Z(n407) );
  XNOR2_X1 U432 ( .A(n406), .B(n408), .ZN(n669) );
  XNOR2_X1 U433 ( .A(n556), .B(n373), .ZN(n751) );
  XNOR2_X1 U434 ( .A(n776), .B(n558), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n409), .B(n520), .ZN(n406) );
  BUF_X1 U436 ( .A(n566), .Z(n408) );
  AND2_X1 U437 ( .A1(n713), .A2(n362), .ZN(n361) );
  NOR2_X1 U438 ( .A1(n366), .A2(n365), .ZN(n364) );
  NAND2_X1 U439 ( .A1(n401), .A2(n400), .ZN(n399) );
  XNOR2_X1 U440 ( .A(n465), .B(n552), .ZN(n776) );
  XNOR2_X1 U441 ( .A(n771), .B(KEYINPUT70), .ZN(n570) );
  XNOR2_X1 U442 ( .A(n529), .B(n418), .ZN(n485) );
  NAND2_X1 U443 ( .A1(n366), .A2(n365), .ZN(n362) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n529) );
  XNOR2_X1 U445 ( .A(n371), .B(n370), .ZN(n555) );
  XNOR2_X1 U446 ( .A(n551), .B(G140), .ZN(n465) );
  XNOR2_X1 U447 ( .A(n356), .B(G107), .ZN(n355) );
  AND2_X1 U448 ( .A1(G214), .A2(n557), .ZN(n558) );
  INV_X1 U449 ( .A(n713), .ZN(n353) );
  XNOR2_X1 U450 ( .A(n392), .B(G116), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n553), .B(G122), .ZN(n371) );
  XNOR2_X1 U452 ( .A(n358), .B(n357), .ZN(n391) );
  XNOR2_X1 U453 ( .A(G101), .B(G110), .ZN(n354) );
  XNOR2_X1 U454 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n370) );
  XOR2_X1 U455 ( .A(G137), .B(KEYINPUT67), .Z(n573) );
  XOR2_X1 U456 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n552) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(KEYINPUT68), .ZN(n358) );
  NOR2_X1 U458 ( .A1(G953), .A2(G237), .ZN(n557) );
  XNOR2_X1 U459 ( .A(G146), .B(G101), .ZN(n517) );
  INV_X1 U460 ( .A(KEYINPUT42), .ZN(n389) );
  NOR2_X1 U461 ( .A1(G902), .A2(n761), .ZN(n585) );
  XNOR2_X2 U462 ( .A(n457), .B(n508), .ZN(n747) );
  XNOR2_X1 U463 ( .A(n367), .B(n649), .ZN(n656) );
  NOR2_X2 U464 ( .A1(n640), .A2(n428), .ZN(n696) );
  INV_X1 U465 ( .A(n570), .ZN(n527) );
  NAND2_X1 U466 ( .A1(n674), .A2(n560), .ZN(n531) );
  NAND2_X1 U467 ( .A1(n674), .A2(n364), .ZN(n363) );
  INV_X1 U468 ( .A(n560), .ZN(n365) );
  XNOR2_X2 U469 ( .A(n644), .B(n533), .ZN(n452) );
  NAND2_X1 U470 ( .A1(n368), .A2(n499), .ZN(n367) );
  XNOR2_X1 U471 ( .A(n369), .B(n501), .ZN(n368) );
  NAND2_X1 U472 ( .A1(n462), .A2(n463), .ZN(n369) );
  NAND2_X1 U473 ( .A1(n503), .A2(n351), .ZN(n388) );
  NAND2_X1 U474 ( .A1(n379), .A2(n389), .ZN(n378) );
  INV_X1 U475 ( .A(n383), .ZN(n379) );
  NAND2_X1 U476 ( .A1(n381), .A2(n389), .ZN(n380) );
  NAND2_X1 U477 ( .A1(n382), .A2(n386), .ZN(n381) );
  INV_X1 U478 ( .A(n640), .ZN(n382) );
  NOR2_X1 U479 ( .A1(n353), .A2(n351), .ZN(n384) );
  INV_X1 U480 ( .A(n503), .ZN(n385) );
  NAND2_X1 U481 ( .A1(n353), .A2(n351), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n396), .A2(n402), .ZN(n394) );
  NAND2_X1 U483 ( .A1(n402), .A2(n398), .ZN(n618) );
  NAND2_X1 U484 ( .A1(n747), .A2(G469), .ZN(n404) );
  BUF_X1 U485 ( .A(n529), .Z(n409) );
  BUF_X2 U486 ( .A(n725), .Z(n410) );
  INV_X1 U487 ( .A(G134), .ZN(n515) );
  XNOR2_X1 U488 ( .A(KEYINPUT4), .B(G131), .ZN(n516) );
  XNOR2_X1 U489 ( .A(n512), .B(n564), .ZN(n589) );
  INV_X1 U490 ( .A(n723), .ZN(n605) );
  INV_X1 U491 ( .A(n456), .ZN(n455) );
  INV_X1 U492 ( .A(KEYINPUT88), .ZN(n451) );
  INV_X1 U493 ( .A(n705), .ZN(n500) );
  INV_X1 U494 ( .A(KEYINPUT65), .ZN(n448) );
  INV_X1 U495 ( .A(KEYINPUT46), .ZN(n501) );
  AND2_X1 U496 ( .A1(n438), .A2(n607), .ZN(n431) );
  XOR2_X1 U497 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n544) );
  XNOR2_X1 U498 ( .A(G107), .B(KEYINPUT9), .ZN(n543) );
  XNOR2_X1 U499 ( .A(n549), .B(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U500 ( .A(G116), .B(G122), .ZN(n542) );
  XOR2_X1 U501 ( .A(G146), .B(G140), .Z(n568) );
  INV_X1 U502 ( .A(n573), .ZN(n565) );
  INV_X1 U503 ( .A(KEYINPUT113), .ZN(n502) );
  XNOR2_X1 U504 ( .A(n637), .B(KEYINPUT39), .ZN(n638) );
  NOR2_X1 U505 ( .A1(G952), .A2(n781), .ZN(n763) );
  NAND2_X1 U506 ( .A1(n471), .A2(n473), .ZN(n472) );
  XNOR2_X1 U507 ( .A(n604), .B(KEYINPUT86), .ZN(n471) );
  NOR2_X1 U508 ( .A1(KEYINPUT87), .A2(n445), .ZN(n444) );
  INV_X1 U509 ( .A(KEYINPUT44), .ZN(n445) );
  NAND2_X1 U510 ( .A1(n440), .A2(n439), .ZN(n438) );
  NOR2_X1 U511 ( .A1(n500), .A2(n415), .ZN(n478) );
  XNOR2_X1 U512 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U513 ( .A(KEYINPUT17), .B(KEYINPUT94), .Z(n525) );
  XNOR2_X1 U514 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n524) );
  XOR2_X1 U515 ( .A(KEYINPUT5), .B(G137), .Z(n518) );
  INV_X1 U516 ( .A(KEYINPUT45), .ZN(n608) );
  NAND2_X1 U517 ( .A1(G234), .A2(G237), .ZN(n534) );
  OR2_X1 U518 ( .A1(G237), .A2(G902), .ZN(n532) );
  INV_X1 U519 ( .A(KEYINPUT38), .ZN(n488) );
  INV_X1 U520 ( .A(KEYINPUT107), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT6), .B(n410), .Z(n641) );
  XOR2_X1 U522 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n530) );
  XOR2_X1 U523 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n575) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(G110), .Z(n572) );
  XNOR2_X1 U525 ( .A(G113), .B(G131), .ZN(n554) );
  NAND2_X1 U526 ( .A1(n622), .A2(n621), .ZN(n461) );
  XNOR2_X1 U527 ( .A(n481), .B(n480), .ZN(n686) );
  INV_X1 U528 ( .A(KEYINPUT99), .ZN(n480) );
  AND2_X1 U529 ( .A1(n622), .A2(n597), .ZN(n598) );
  NOR2_X1 U530 ( .A1(n589), .A2(n641), .ZN(n604) );
  XNOR2_X1 U531 ( .A(n506), .B(n504), .ZN(n756) );
  XNOR2_X1 U532 ( .A(n505), .B(n547), .ZN(n504) );
  XNOR2_X1 U533 ( .A(n546), .B(n419), .ZN(n506) );
  XNOR2_X1 U534 ( .A(n570), .B(n569), .ZN(n508) );
  XNOR2_X1 U535 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U536 ( .A1(n657), .A2(n697), .ZN(n464) );
  INV_X1 U537 ( .A(n730), .ZN(n454) );
  XNOR2_X1 U538 ( .A(KEYINPUT106), .B(n588), .ZN(n793) );
  INV_X1 U539 ( .A(n763), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n745), .B(n479), .ZN(G75) );
  XNOR2_X1 U541 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n479) );
  INV_X1 U542 ( .A(n472), .ZN(n683) );
  AND2_X1 U543 ( .A1(n792), .A2(n660), .ZN(n411) );
  AND2_X1 U544 ( .A1(n792), .A2(n423), .ZN(n412) );
  AND2_X1 U545 ( .A1(n435), .A2(n667), .ZN(n413) );
  AND2_X1 U546 ( .A1(G210), .A2(n532), .ZN(n414) );
  AND2_X1 U547 ( .A1(n633), .A2(n696), .ZN(n415) );
  XNOR2_X1 U548 ( .A(n626), .B(KEYINPUT77), .ZN(n416) );
  AND2_X1 U549 ( .A1(n667), .A2(G475), .ZN(n417) );
  XOR2_X1 U550 ( .A(n530), .B(G122), .Z(n418) );
  AND2_X1 U551 ( .A1(G217), .A2(n578), .ZN(n419) );
  AND2_X1 U552 ( .A1(n450), .A2(KEYINPUT87), .ZN(n420) );
  XNOR2_X1 U553 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n421) );
  XOR2_X1 U554 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n422) );
  XOR2_X1 U555 ( .A(G902), .B(KEYINPUT15), .Z(n660) );
  AND2_X1 U556 ( .A1(n660), .A2(n497), .ZN(n423) );
  XOR2_X1 U557 ( .A(n608), .B(KEYINPUT83), .Z(n424) );
  XOR2_X1 U558 ( .A(n671), .B(n670), .Z(n425) );
  INV_X1 U559 ( .A(KEYINPUT87), .ZN(n607) );
  INV_X1 U560 ( .A(KEYINPUT82), .ZN(n497) );
  NAND2_X1 U561 ( .A1(n426), .A2(n454), .ZN(n453) );
  NAND2_X1 U562 ( .A1(n563), .A2(n426), .ZN(n512) );
  XNOR2_X2 U563 ( .A(n541), .B(n540), .ZN(n426) );
  INV_X1 U564 ( .A(n492), .ZN(n427) );
  BUF_X1 U565 ( .A(n452), .Z(n428) );
  XNOR2_X1 U566 ( .A(n531), .B(n414), .ZN(n429) );
  AND2_X1 U567 ( .A1(n793), .A2(n788), .ZN(n430) );
  NAND2_X1 U568 ( .A1(n441), .A2(n431), .ZN(n458) );
  NAND2_X1 U569 ( .A1(n441), .A2(n438), .ZN(n432) );
  NAND2_X1 U570 ( .A1(n493), .A2(n491), .ZN(n433) );
  NAND2_X1 U571 ( .A1(n493), .A2(n491), .ZN(n662) );
  AND2_X2 U572 ( .A1(n496), .A2(n494), .ZN(n493) );
  XNOR2_X1 U573 ( .A(n600), .B(n460), .ZN(n592) );
  BUF_X1 U574 ( .A(n644), .Z(n434) );
  XNOR2_X1 U575 ( .A(n593), .B(KEYINPUT33), .ZN(n706) );
  INV_X1 U576 ( .A(n410), .ZN(n597) );
  AND2_X1 U577 ( .A1(n667), .A2(G210), .ZN(n510) );
  NOR2_X1 U578 ( .A1(n719), .A2(n723), .ZN(n473) );
  NAND2_X1 U579 ( .A1(n433), .A2(n661), .ZN(n435) );
  NAND2_X1 U580 ( .A1(n662), .A2(n661), .ZN(n668) );
  AND2_X1 U581 ( .A1(n436), .A2(n447), .ZN(n446) );
  NAND2_X1 U582 ( .A1(n437), .A2(n430), .ZN(n436) );
  XNOR2_X1 U583 ( .A(n596), .B(n448), .ZN(n437) );
  INV_X1 U584 ( .A(n469), .ZN(n439) );
  NOR2_X1 U585 ( .A1(n468), .A2(n451), .ZN(n440) );
  AND2_X2 U586 ( .A1(n442), .A2(n443), .ZN(n441) );
  NAND2_X1 U587 ( .A1(n468), .A2(n451), .ZN(n442) );
  NAND2_X1 U588 ( .A1(n469), .A2(n451), .ZN(n443) );
  NAND2_X1 U589 ( .A1(n606), .A2(KEYINPUT44), .ZN(n450) );
  NAND2_X1 U590 ( .A1(n606), .A2(n444), .ZN(n447) );
  AND2_X2 U591 ( .A1(n449), .A2(n446), .ZN(n459) );
  NAND2_X1 U592 ( .A1(n432), .A2(n420), .ZN(n449) );
  NOR2_X2 U593 ( .A1(n452), .A2(n539), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n455), .A2(n686), .ZN(n601) );
  AND2_X1 U595 ( .A1(n456), .A2(n691), .ZN(n703) );
  AND2_X1 U596 ( .A1(n456), .A2(n697), .ZN(n701) );
  INV_X1 U597 ( .A(n667), .ZN(n740) );
  OR2_X2 U598 ( .A1(n764), .A2(n666), .ZN(n667) );
  XNOR2_X2 U599 ( .A(n566), .B(n565), .ZN(n457) );
  XNOR2_X1 U600 ( .A(n407), .B(n776), .ZN(n780) );
  NAND2_X2 U601 ( .A1(n459), .A2(n458), .ZN(n474) );
  XNOR2_X1 U602 ( .A(n461), .B(KEYINPUT75), .ZN(n625) );
  AND2_X1 U603 ( .A1(n720), .A2(n618), .ZN(n622) );
  INV_X1 U604 ( .A(n791), .ZN(n462) );
  INV_X1 U605 ( .A(n785), .ZN(n463) );
  XNOR2_X2 U606 ( .A(n466), .B(G125), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n467), .A2(n631), .ZN(n470) );
  XNOR2_X1 U608 ( .A(n601), .B(KEYINPUT100), .ZN(n467) );
  XNOR2_X2 U609 ( .A(n482), .B(KEYINPUT35), .ZN(n787) );
  NAND2_X1 U610 ( .A1(n470), .A2(n472), .ZN(n469) );
  XNOR2_X2 U611 ( .A(n474), .B(n424), .ZN(n764) );
  BUF_X1 U612 ( .A(n686), .Z(n475) );
  NAND2_X1 U613 ( .A1(n599), .A2(n598), .ZN(n481) );
  XNOR2_X1 U614 ( .A(n672), .B(n425), .ZN(n477) );
  NOR2_X1 U615 ( .A1(n679), .A2(n763), .ZN(n682) );
  NOR2_X1 U616 ( .A1(n754), .A2(n763), .ZN(n755) );
  NAND2_X1 U617 ( .A1(n477), .A2(n476), .ZN(n673) );
  NOR2_X1 U618 ( .A1(KEYINPUT2), .A2(n498), .ZN(n739) );
  NOR2_X1 U619 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U620 ( .A1(n659), .A2(n792), .ZN(n779) );
  INV_X1 U621 ( .A(n764), .ZN(n492) );
  XNOR2_X1 U622 ( .A(n594), .B(n421), .ZN(n483) );
  NAND2_X1 U623 ( .A1(n483), .A2(n416), .ZN(n482) );
  INV_X1 U624 ( .A(n485), .ZN(n770) );
  XNOR2_X1 U625 ( .A(n487), .B(n526), .ZN(n486) );
  XNOR2_X1 U626 ( .A(n551), .B(n523), .ZN(n487) );
  INV_X1 U627 ( .A(n429), .ZN(n653) );
  XNOR2_X1 U628 ( .A(n653), .B(n488), .ZN(n635) );
  NAND2_X1 U629 ( .A1(n627), .A2(n429), .ZN(n695) );
  NAND2_X1 U630 ( .A1(n659), .A2(n412), .ZN(n490) );
  NAND2_X1 U631 ( .A1(n489), .A2(KEYINPUT82), .ZN(n494) );
  NAND2_X1 U632 ( .A1(n659), .A2(n411), .ZN(n489) );
  INV_X1 U633 ( .A(n779), .ZN(n495) );
  NAND2_X1 U634 ( .A1(n764), .A2(KEYINPUT82), .ZN(n496) );
  XNOR2_X2 U635 ( .A(n545), .B(n516), .ZN(n566) );
  XNOR2_X2 U636 ( .A(n507), .B(G143), .ZN(n528) );
  NAND2_X1 U637 ( .A1(n668), .A2(n510), .ZN(n678) );
  NAND2_X1 U638 ( .A1(n668), .A2(n417), .ZN(n752) );
  NAND2_X1 U639 ( .A1(n435), .A2(n511), .ZN(n672) );
  AND2_X1 U640 ( .A1(n667), .A2(G472), .ZN(n511) );
  NAND2_X1 U641 ( .A1(n413), .A2(G217), .ZN(n760) );
  NAND2_X1 U642 ( .A1(n413), .A2(G478), .ZN(n757) );
  NAND2_X1 U643 ( .A1(n413), .A2(G469), .ZN(n749) );
  AND2_X1 U644 ( .A1(G221), .A2(n578), .ZN(n513) );
  AND2_X1 U645 ( .A1(n557), .A2(G210), .ZN(n514) );
  INV_X1 U646 ( .A(KEYINPUT91), .ZN(n521) );
  XNOR2_X1 U647 ( .A(n519), .B(n514), .ZN(n520) );
  BUF_X1 U648 ( .A(n706), .Z(n717) );
  INV_X1 U649 ( .A(KEYINPUT85), .ZN(n637) );
  XNOR2_X1 U650 ( .A(KEYINPUT64), .B(KEYINPUT22), .ZN(n564) );
  XNOR2_X1 U651 ( .A(n776), .B(n513), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n580), .B(n579), .ZN(n761) );
  XNOR2_X1 U653 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U654 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U655 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U656 ( .A(n660), .ZN(n560) );
  NAND2_X1 U657 ( .A1(G224), .A2(n781), .ZN(n522) );
  XNOR2_X1 U658 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U659 ( .A1(G214), .A2(n532), .ZN(n713) );
  XOR2_X1 U660 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n533) );
  XNOR2_X1 U661 ( .A(KEYINPUT14), .B(n534), .ZN(n536) );
  NAND2_X1 U662 ( .A1(G952), .A2(n536), .ZN(n738) );
  NOR2_X1 U663 ( .A1(G953), .A2(n738), .ZN(n535) );
  XOR2_X1 U664 ( .A(KEYINPUT95), .B(n535), .Z(n612) );
  AND2_X1 U665 ( .A1(G953), .A2(n536), .ZN(n537) );
  NAND2_X1 U666 ( .A1(G902), .A2(n537), .ZN(n609) );
  NOR2_X1 U667 ( .A1(n609), .A2(G898), .ZN(n538) );
  NOR2_X1 U668 ( .A1(n612), .A2(n538), .ZN(n539) );
  XNOR2_X1 U669 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U670 ( .A(n542), .B(KEYINPUT101), .ZN(n549) );
  XNOR2_X1 U671 ( .A(n544), .B(n543), .ZN(n547) );
  XNOR2_X1 U672 ( .A(n545), .B(KEYINPUT103), .ZN(n546) );
  NAND2_X1 U673 ( .A1(G234), .A2(n781), .ZN(n548) );
  XOR2_X1 U674 ( .A(KEYINPUT8), .B(n548), .Z(n578) );
  NOR2_X1 U675 ( .A1(G902), .A2(n756), .ZN(n550) );
  XOR2_X1 U676 ( .A(G478), .B(n550), .Z(n595) );
  XNOR2_X1 U677 ( .A(n555), .B(n554), .ZN(n556) );
  NOR2_X1 U678 ( .A1(n595), .A2(n602), .ZN(n559) );
  NAND2_X1 U679 ( .A1(n560), .A2(G234), .ZN(n561) );
  XNOR2_X1 U680 ( .A(n561), .B(KEYINPUT20), .ZN(n581) );
  NAND2_X1 U681 ( .A1(n581), .A2(G221), .ZN(n562) );
  XNOR2_X1 U682 ( .A(KEYINPUT21), .B(n562), .ZN(n722) );
  NOR2_X1 U683 ( .A1(n711), .A2(n722), .ZN(n563) );
  NOR2_X1 U684 ( .A1(n589), .A2(n410), .ZN(n587) );
  NAND2_X1 U685 ( .A1(G227), .A2(n781), .ZN(n567) );
  XNOR2_X1 U686 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U687 ( .A(n572), .B(n571), .ZN(n577) );
  XNOR2_X1 U688 ( .A(n573), .B(KEYINPUT81), .ZN(n574) );
  XNOR2_X1 U689 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U690 ( .A(n577), .B(n576), .Z(n580) );
  XOR2_X1 U691 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n583) );
  NAND2_X1 U692 ( .A1(G217), .A2(n581), .ZN(n582) );
  XNOR2_X1 U693 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X2 U694 ( .A(n585), .B(n584), .ZN(n723) );
  NOR2_X1 U695 ( .A1(n719), .A2(n605), .ZN(n586) );
  NAND2_X1 U696 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U697 ( .A(KEYINPUT93), .B(n719), .Z(n648) );
  AND2_X1 U698 ( .A1(n723), .A2(n648), .ZN(n590) );
  NAND2_X1 U699 ( .A1(n604), .A2(n590), .ZN(n591) );
  NAND2_X1 U700 ( .A1(n793), .A2(n788), .ZN(n606) );
  NAND2_X1 U701 ( .A1(n592), .A2(n641), .ZN(n593) );
  NAND2_X1 U702 ( .A1(n706), .A2(n599), .ZN(n594) );
  NAND2_X1 U703 ( .A1(n602), .A2(n595), .ZN(n626) );
  NOR2_X1 U704 ( .A1(n787), .A2(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U705 ( .A1(n410), .A2(n600), .ZN(n730) );
  INV_X1 U706 ( .A(n602), .ZN(n603) );
  INV_X1 U707 ( .A(n697), .ZN(n699) );
  NAND2_X1 U708 ( .A1(n595), .A2(n603), .ZN(n702) );
  NAND2_X1 U709 ( .A1(n699), .A2(n702), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n609), .B(KEYINPUT108), .ZN(n610) );
  NOR2_X1 U711 ( .A1(G900), .A2(n610), .ZN(n611) );
  XNOR2_X1 U712 ( .A(n611), .B(KEYINPUT109), .ZN(n614) );
  INV_X1 U713 ( .A(n612), .ZN(n613) );
  NAND2_X1 U714 ( .A1(n614), .A2(n613), .ZN(n621) );
  NAND2_X1 U715 ( .A1(n723), .A2(n621), .ZN(n615) );
  NAND2_X1 U716 ( .A1(n410), .A2(n643), .ZN(n616) );
  XNOR2_X1 U717 ( .A(KEYINPUT111), .B(n617), .ZN(n619) );
  NAND2_X1 U718 ( .A1(n619), .A2(n618), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n631), .A2(n696), .ZN(n620) );
  NAND2_X1 U720 ( .A1(n620), .A2(KEYINPUT47), .ZN(n629) );
  NAND2_X1 U721 ( .A1(n410), .A2(n713), .ZN(n623) );
  XOR2_X1 U722 ( .A(KEYINPUT30), .B(n623), .Z(n624) );
  NAND2_X1 U723 ( .A1(n625), .A2(n624), .ZN(n636) );
  NOR2_X1 U724 ( .A1(n636), .A2(n626), .ZN(n627) );
  XNOR2_X1 U725 ( .A(KEYINPUT80), .B(n695), .ZN(n628) );
  NAND2_X1 U726 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U727 ( .A(n630), .B(KEYINPUT79), .ZN(n634) );
  INV_X1 U728 ( .A(n631), .ZN(n710) );
  NOR2_X1 U729 ( .A1(KEYINPUT47), .A2(n710), .ZN(n632) );
  XOR2_X1 U730 ( .A(KEYINPUT73), .B(n632), .Z(n633) );
  XNOR2_X1 U731 ( .A(n635), .B(KEYINPUT74), .ZN(n709) );
  OR2_X1 U732 ( .A1(n636), .A2(n709), .ZN(n639) );
  AND2_X1 U733 ( .A1(n697), .A2(n641), .ZN(n642) );
  NAND2_X1 U734 ( .A1(n643), .A2(n642), .ZN(n650) );
  NOR2_X1 U735 ( .A1(n650), .A2(n434), .ZN(n646) );
  XOR2_X1 U736 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n645) );
  XNOR2_X1 U737 ( .A(n646), .B(n645), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n705) );
  XOR2_X1 U739 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n649) );
  NOR2_X1 U740 ( .A1(n719), .A2(n650), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n651), .A2(n713), .ZN(n652) );
  XNOR2_X1 U742 ( .A(n652), .B(KEYINPUT43), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U744 ( .A(KEYINPUT110), .B(n655), .ZN(n790) );
  NAND2_X1 U745 ( .A1(n656), .A2(n790), .ZN(n665) );
  INV_X1 U746 ( .A(n702), .ZN(n691) );
  NAND2_X1 U747 ( .A1(n691), .A2(n657), .ZN(n658) );
  XNOR2_X1 U748 ( .A(n658), .B(KEYINPUT114), .ZN(n792) );
  NAND2_X1 U749 ( .A1(KEYINPUT2), .A2(n660), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n792), .A2(KEYINPUT2), .ZN(n663) );
  XNOR2_X1 U751 ( .A(KEYINPUT78), .B(n663), .ZN(n664) );
  XNOR2_X1 U752 ( .A(n669), .B(KEYINPUT115), .ZN(n671) );
  XOR2_X1 U753 ( .A(KEYINPUT62), .B(KEYINPUT92), .Z(n670) );
  XNOR2_X1 U754 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U755 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT122), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n678), .B(n677), .ZN(n679) );
  INV_X1 U758 ( .A(KEYINPUT123), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n680), .B(KEYINPUT56), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n682), .B(n681), .ZN(G51) );
  XOR2_X1 U761 ( .A(n683), .B(G101), .Z(n684) );
  XNOR2_X1 U762 ( .A(KEYINPUT116), .B(n684), .ZN(G3) );
  NOR2_X1 U763 ( .A1(n699), .A2(n475), .ZN(n685) );
  XOR2_X1 U764 ( .A(G104), .B(n685), .Z(G6) );
  NOR2_X1 U765 ( .A1(n475), .A2(n702), .ZN(n690) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n688) );
  XNOR2_X1 U767 ( .A(G107), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U768 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U769 ( .A(n690), .B(n689), .ZN(G9) );
  XOR2_X1 U770 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n693) );
  NAND2_X1 U771 ( .A1(n691), .A2(n696), .ZN(n692) );
  XNOR2_X1 U772 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U773 ( .A(G128), .B(n694), .ZN(G30) );
  XNOR2_X1 U774 ( .A(G143), .B(n695), .ZN(G45) );
  NAND2_X1 U775 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U776 ( .A(G146), .B(n698), .ZN(G48) );
  XNOR2_X1 U777 ( .A(G113), .B(KEYINPUT119), .ZN(n700) );
  XNOR2_X1 U778 ( .A(n701), .B(n700), .ZN(G15) );
  XOR2_X1 U779 ( .A(G116), .B(n703), .Z(G18) );
  XOR2_X1 U780 ( .A(G125), .B(KEYINPUT37), .Z(n704) );
  XNOR2_X1 U781 ( .A(n705), .B(n704), .ZN(G27) );
  INV_X1 U782 ( .A(n717), .ZN(n707) );
  NOR2_X1 U783 ( .A1(n733), .A2(n707), .ZN(n708) );
  NOR2_X1 U784 ( .A1(G953), .A2(n708), .ZN(n744) );
  OR2_X1 U785 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U787 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U788 ( .A1(n503), .A2(n715), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U790 ( .A(KEYINPUT120), .B(n718), .Z(n735) );
  NOR2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U792 ( .A(KEYINPUT50), .B(n721), .Z(n728) );
  NAND2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U794 ( .A(n724), .B(KEYINPUT49), .ZN(n726) );
  NOR2_X1 U795 ( .A1(n726), .A2(n410), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U798 ( .A(KEYINPUT51), .B(n731), .ZN(n732) );
  NOR2_X1 U799 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U800 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U801 ( .A(n736), .B(KEYINPUT52), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n738), .A2(n737), .ZN(n742) );
  NOR2_X1 U803 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U804 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  NOR2_X1 U806 ( .A1(n763), .A2(n750), .ZN(G54) );
  XOR2_X1 U807 ( .A(n751), .B(KEYINPUT59), .Z(n753) );
  XNOR2_X1 U808 ( .A(n752), .B(n753), .ZN(n754) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U810 ( .A(n756), .B(KEYINPUT124), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n763), .A2(n759), .ZN(G63) );
  XNOR2_X1 U813 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n763), .A2(n762), .ZN(G66) );
  NOR2_X1 U815 ( .A1(G953), .A2(n427), .ZN(n765) );
  XNOR2_X1 U816 ( .A(KEYINPUT125), .B(n765), .ZN(n769) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U820 ( .A1(n769), .A2(n768), .ZN(n775) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n773) );
  NOR2_X1 U822 ( .A1(n781), .A2(G898), .ZN(n772) );
  NOR2_X1 U823 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(G69) );
  XNOR2_X1 U825 ( .A(G227), .B(n780), .ZN(n777) );
  NAND2_X1 U826 ( .A1(G900), .A2(n777), .ZN(n778) );
  NAND2_X1 U827 ( .A1(n778), .A2(G953), .ZN(n784) );
  XNOR2_X1 U828 ( .A(n780), .B(n779), .ZN(n782) );
  NAND2_X1 U829 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(G72) );
  XNOR2_X1 U831 ( .A(n785), .B(G131), .ZN(n786) );
  XNOR2_X1 U832 ( .A(n786), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U833 ( .A(n787), .B(G122), .Z(G24) );
  XNOR2_X1 U834 ( .A(G119), .B(n788), .ZN(n789) );
  XNOR2_X1 U835 ( .A(n789), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U836 ( .A(G140), .B(n790), .ZN(G42) );
  XOR2_X1 U837 ( .A(G137), .B(n791), .Z(G39) );
  XNOR2_X1 U838 ( .A(G134), .B(n792), .ZN(G36) );
  XNOR2_X1 U839 ( .A(G110), .B(n793), .ZN(G12) );
endmodule

