//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g028(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n455), .A2(new_n451), .B1(new_n459), .B2(new_n456), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT69), .B1(new_n463), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n475), .A2(KEYINPUT70), .A3(G101), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n471), .B2(new_n474), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n470), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n473), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(G160));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n473), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n473), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n486), .A2(new_n504), .A3(G138), .A4(new_n473), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n512), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n511), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  OAI211_X1 g102(.A(G543), .B(new_n519), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n528), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT73), .A3(G50), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n522), .A2(new_n524), .A3(new_n530), .A4(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n520), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n539), .B(new_n543), .C1(new_n528), .C2(new_n540), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n538), .B1(new_n542), .B2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n521), .A2(G90), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n511), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n531), .A2(G52), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n514), .A2(new_n516), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(new_n526), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(new_n557));
  AOI22_X1  g132(.A1(new_n521), .A2(G81), .B1(G43), .B2(new_n531), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n553), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT77), .ZN(new_n570));
  XOR2_X1   g145(.A(KEYINPUT78), .B(G65), .Z(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n507), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n518), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n575), .A2(G91), .A3(new_n517), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n528), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n575), .A2(new_n581), .A3(G53), .A4(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT79), .B1(new_n578), .B2(new_n583), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G299));
  AND2_X1   g163(.A1(G168), .A2(KEYINPUT80), .ZN(new_n589));
  NOR2_X1   g164(.A1(G168), .A2(KEYINPUT80), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G286));
  OAI21_X1  g167(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G49), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n528), .B2(new_n594), .C1(new_n520), .C2(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n553), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(new_n526), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n602), .A3(new_n526), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n601), .A2(new_n603), .B1(new_n531), .B2(G48), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n575), .A2(G86), .A3(new_n517), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT82), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n575), .A2(new_n607), .A3(G86), .A4(new_n517), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n604), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(G72), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G60), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n553), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n531), .A2(G47), .B1(new_n526), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n521), .A2(G85), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT10), .B1(new_n520), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n575), .A2(new_n620), .A3(G92), .A4(new_n517), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT77), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT77), .B1(new_n514), .B2(new_n516), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G66), .ZN(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n507), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n531), .A2(G54), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n617), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n617), .B1(new_n630), .B2(G868), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n591), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n587), .B(KEYINPUT84), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(G868), .B2(new_n636), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(G868), .B2(new_n636), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n559), .A2(new_n633), .ZN(new_n641));
  INV_X1    g216(.A(new_n630), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n642), .A2(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n643), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n475), .A2(new_n486), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  OR2_X1    g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n651));
  INV_X1    g226(.A(G135), .ZN(new_n652));
  INV_X1    g227(.A(G123), .ZN(new_n653));
  OAI221_X1 g228(.A(new_n651), .B1(new_n490), .B2(new_n652), .C1(new_n653), .C2(new_n487), .ZN(new_n654));
  INV_X1    g229(.A(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT15), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(G2435), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(G2435), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(G14), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT17), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n655), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(G2100), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT87), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(KEYINPUT87), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n687), .A2(new_n689), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n698), .A2(new_n699), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n696), .A2(new_n691), .A3(new_n700), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(new_n699), .C2(new_n698), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT88), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(G1981), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(G1991), .B(G1996), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n706), .B(new_n711), .ZN(G229));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G107), .B2(new_n473), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT91), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n488), .A2(G119), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n491), .A2(G131), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(G29), .ZN(new_n722));
  MUX2_X1   g297(.A(new_n714), .B(new_n722), .S(KEYINPUT90), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n723), .B(new_n725), .Z(new_n726));
  MUX2_X1   g301(.A(G24), .B(G290), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G23), .ZN(new_n730));
  INV_X1    g305(.A(G288), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT33), .B(G1976), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n735), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G1971), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G1971), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n735), .A2(G6), .ZN(new_n742));
  INV_X1    g317(.A(G305), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n735), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT32), .B(G1981), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT34), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n747), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n749), .A2(new_n740), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n729), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT36), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(new_n729), .C1(new_n748), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n713), .A2(G35), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n495), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT31), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n760), .A2(G2090), .B1(new_n761), .B2(G11), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(G11), .ZN(new_n763));
  NOR2_X1   g338(.A1(G164), .A2(new_n713), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G27), .B2(new_n713), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G2078), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(G2078), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT27), .B(G1996), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT97), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n488), .A2(G129), .B1(G105), .B2(new_n475), .ZN(new_n771));
  INV_X1    g346(.A(G141), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n490), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G32), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n767), .B(new_n768), .C1(new_n770), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n735), .A2(KEYINPUT23), .A3(G20), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n783));
  INV_X1    g358(.A(G20), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G16), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n785), .C1(new_n587), .C2(new_n735), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n760), .A2(G2090), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT98), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  NAND2_X1  g367(.A1(G168), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G16), .B2(G21), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n735), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n630), .B2(new_n735), .ZN(new_n798));
  INV_X1    g373(.A(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n788), .A2(new_n795), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT30), .B(G28), .Z(new_n802));
  OAI22_X1  g377(.A1(new_n780), .A2(new_n770), .B1(G29), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT25), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G139), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n490), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT94), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n809), .A2(new_n810), .B1(new_n473), .B2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G33), .B(new_n812), .S(G29), .Z(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G2072), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n735), .A2(G5), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G171), .B2(new_n735), .ZN(new_n816));
  INV_X1    g391(.A(G1961), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n735), .A2(G19), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n560), .B2(new_n735), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1341), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n801), .A2(new_n803), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n756), .A2(new_n763), .A3(new_n781), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT28), .ZN(new_n825));
  INV_X1    g400(.A(G26), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G29), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(G29), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n488), .A2(G128), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n491), .A2(G140), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n473), .A2(G116), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n828), .B1(new_n833), .B2(G29), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n827), .B1(new_n834), .B2(new_n825), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n654), .A2(new_n713), .ZN(new_n837));
  OR2_X1    g412(.A1(KEYINPUT24), .A2(G34), .ZN(new_n838));
  NAND2_X1  g413(.A1(KEYINPUT24), .A2(G34), .ZN(new_n839));
  AOI21_X1  g414(.A(G29), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G160), .B2(G29), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT95), .B(G2084), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n824), .A2(new_n836), .A3(new_n837), .A4(new_n843), .ZN(G311));
  AND4_X1   g419(.A1(new_n756), .A2(new_n763), .A3(new_n781), .A4(new_n823), .ZN(new_n845));
  INV_X1    g420(.A(new_n836), .ZN(new_n846));
  INV_X1    g421(.A(new_n837), .ZN(new_n847));
  INV_X1    g422(.A(new_n843), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(G150));
  XNOR2_X1  g424(.A(KEYINPUT99), .B(G93), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n521), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n511), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n531), .A2(G55), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n559), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n630), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n857), .B1(new_n863), .B2(G860), .ZN(G145));
  NAND2_X1  g439(.A1(new_n503), .A2(new_n505), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n497), .A2(new_n500), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n812), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n833), .ZN(new_n869));
  INV_X1    g444(.A(new_n778), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  AOI22_X1  g448(.A1(G130), .A2(new_n488), .B1(new_n491), .B2(G142), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n473), .A2(G118), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT100), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n721), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n647), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n879), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n647), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n881), .B2(new_n885), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n872), .B(new_n873), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n873), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n891), .A2(new_n871), .B1(new_n886), .B2(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G160), .B(new_n495), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n654), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n897), .A2(new_n902), .A3(new_n899), .A4(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(G395));
  XOR2_X1   g479(.A(new_n859), .B(new_n643), .Z(new_n905));
  OAI21_X1  g480(.A(new_n642), .B1(new_n585), .B2(new_n586), .ZN(new_n906));
  INV_X1    g481(.A(new_n586), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n630), .A3(new_n584), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n905), .A2(KEYINPUT103), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(new_n905), .B2(new_n909), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n906), .B2(new_n908), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n905), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G166), .B(G305), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(G288), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G305), .B(G303), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(new_n918), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n920), .A2(new_n922), .A3(KEYINPUT42), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n918), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n929), .B2(KEYINPUT42), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n916), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n916), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g509(.A(new_n933), .B1(G868), .B2(new_n858), .ZN(G331));
  INV_X1    g510(.A(new_n909), .ZN(new_n936));
  OAI21_X1  g511(.A(G171), .B1(new_n589), .B2(new_n590), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT105), .B1(G168), .B2(G301), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(G171), .C1(new_n589), .C2(new_n590), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n859), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n859), .B1(new_n940), .B2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n859), .ZN(new_n947));
  OR2_X1    g522(.A1(G168), .A2(KEYINPUT80), .ZN(new_n948));
  NAND2_X1  g523(.A1(G168), .A2(KEYINPUT80), .ZN(new_n949));
  AOI21_X1  g524(.A(G301), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n938), .ZN(new_n951));
  INV_X1    g526(.A(new_n942), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n914), .A2(new_n953), .A3(new_n943), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n946), .A2(new_n954), .A3(new_n929), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n929), .B1(new_n946), .B2(new_n954), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(new_n956), .A3(G37), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n946), .A2(new_n954), .ZN(new_n960));
  INV_X1    g535(.A(new_n929), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n946), .A2(new_n954), .A3(new_n929), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n898), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n946), .A2(new_n954), .A3(KEYINPUT106), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(new_n898), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n956), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n958), .A3(new_n970), .A4(new_n963), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n966), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n963), .A2(new_n967), .A3(new_n898), .ZN(new_n973));
  AOI211_X1 g548(.A(KEYINPUT106), .B(new_n929), .C1(new_n946), .C2(new_n954), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n962), .A2(new_n958), .A3(new_n898), .A4(new_n963), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(G397));
  XNOR2_X1  g555(.A(new_n478), .B(KEYINPUT70), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n481), .B(KEYINPUT68), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(G40), .A3(new_n470), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G164), .B2(G1384), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n778), .B(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2067), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n833), .B(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n721), .A2(new_n725), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n833), .A2(G2067), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n986), .B1(new_n992), .B2(new_n870), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n986), .A2(KEYINPUT46), .A3(new_n988), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n987), .B2(G1996), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT47), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n721), .A2(new_n725), .ZN(new_n1004));
  INV_X1    g579(.A(new_n994), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n993), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n986), .ZN(new_n1007));
  OR2_X1    g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n987), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n997), .B(new_n1003), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n480), .A2(new_n1013), .A3(new_n483), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n985), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1971), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1020));
  AOI211_X1 g595(.A(KEYINPUT50), .B(G1384), .C1(new_n865), .C2(new_n866), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n867), .A2(new_n1015), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT108), .A3(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1014), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1026), .B2(G2090), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(G166), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(new_n1032), .A3(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n983), .A2(new_n1024), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(G288), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n601), .A2(new_n603), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n531), .A2(G48), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n609), .A2(new_n1039), .A3(new_n708), .A4(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n599), .A2(new_n602), .A3(new_n526), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n602), .B1(new_n599), .B2(new_n526), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(new_n605), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G1981), .ZN(new_n1045));
  OR2_X1    g620(.A1(KEYINPUT109), .A2(KEYINPUT49), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(KEYINPUT109), .A2(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1041), .A2(new_n1045), .A3(KEYINPUT109), .A4(KEYINPUT49), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1035), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1035), .B(new_n1052), .C1(new_n1036), .C2(G288), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1033), .A2(new_n1038), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1032), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n867), .A2(new_n1056), .A3(new_n1057), .A4(new_n1015), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1058), .A2(new_n1020), .ZN(new_n1059));
  INV_X1    g634(.A(G2090), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT111), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1014), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1019), .A3(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT112), .B1(new_n1062), .B2(new_n1019), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1055), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1020), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n865), .B2(new_n866), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1056), .B1(new_n1071), .B2(new_n1057), .ZN(new_n1072));
  NOR4_X1   g647(.A1(new_n1070), .A2(new_n1072), .A3(G2090), .A4(new_n983), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(KEYINPUT45), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n983), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1971), .B1(new_n1075), .B2(new_n1016), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1069), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(new_n1063), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT113), .A3(new_n1055), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1054), .B1(new_n1068), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1026), .A2(new_n817), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1017), .B2(G2078), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT123), .B1(new_n1074), .B2(new_n983), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n484), .A2(new_n985), .A3(new_n1085), .A4(G40), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1082), .A2(G2078), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1016), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1092), .A3(KEYINPUT45), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1075), .A2(new_n1087), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1081), .A2(new_n1083), .A3(G301), .A4(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(KEYINPUT54), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1090), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n1102), .B2(new_n1094), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1089), .A2(G171), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1091), .A2(new_n1014), .A3(new_n985), .A4(new_n1093), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n792), .ZN(new_n1108));
  INV_X1    g683(.A(G2084), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1023), .A2(new_n1109), .A3(new_n1014), .A4(new_n1025), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(G168), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1106), .B1(new_n1111), .B2(G8), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(G168), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1111), .C1(new_n1114), .C2(new_n1106), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1080), .A2(new_n1100), .A3(new_n1105), .A4(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1061), .A2(new_n1014), .A3(new_n1020), .A4(new_n1058), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n787), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1014), .A2(new_n985), .A3(new_n1016), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n578), .B2(new_n583), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n625), .A2(new_n571), .B1(G78), .B2(G543), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n576), .C1(new_n1127), .C2(new_n507), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n574), .B2(new_n577), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT57), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n580), .A2(new_n1131), .A3(new_n582), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n580), .B2(new_n582), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g709(.A(KEYINPUT117), .B(new_n1125), .C1(new_n1130), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1134), .A3(new_n1124), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1125), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1123), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1123), .B(KEYINPUT119), .C1(new_n1135), .C2(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1026), .A2(new_n799), .B1(new_n990), .B2(new_n1034), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n642), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1138), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n787), .A2(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT118), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1149), .A2(new_n1151), .A3(new_n1154), .A4(new_n1150), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1147), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1120), .A2(new_n988), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(G1341), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n983), .B2(new_n1024), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n559), .B(new_n1157), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g738(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n560), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1165), .B2(new_n1157), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1152), .A2(KEYINPUT61), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1145), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1153), .A2(new_n1141), .A3(new_n1155), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n630), .B1(new_n1146), .B2(KEYINPUT60), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT122), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1174), .B(new_n630), .C1(new_n1146), .C2(KEYINPUT60), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1173), .A2(KEYINPUT60), .A3(new_n1146), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1146), .A2(KEYINPUT60), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1168), .A2(new_n1171), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1117), .B1(new_n1156), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1113), .A2(new_n1115), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1054), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1079), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT113), .B1(new_n1078), .B2(new_n1055), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1184), .B(new_n1185), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1114), .A2(new_n1106), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1111), .A2(G8), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1112), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1103), .B1(new_n1192), .B2(new_n1183), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1182), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1103), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n1116), .B2(KEYINPUT62), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1080), .A2(new_n1196), .A3(KEYINPUT125), .A4(new_n1184), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1051), .A2(new_n1036), .A3(new_n731), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1199), .A2(KEYINPUT110), .A3(new_n1041), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT110), .B1(new_n1199), .B2(new_n1041), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1038), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1032), .B1(new_n1027), .B2(G8), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1205), .A2(G8), .A3(new_n591), .ZN(new_n1206));
  OR3_X1    g781(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1202), .A2(new_n1035), .B1(KEYINPUT63), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1033), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1206), .A2(KEYINPUT63), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1208), .B1(new_n1212), .B2(new_n1203), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1181), .A2(new_n1198), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1006), .B1(G1986), .B2(G290), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n987), .B1(new_n1215), .B2(new_n1008), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1012), .B1(new_n1214), .B2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g792(.A1(G229), .A2(new_n460), .ZN(new_n1219));
  AOI21_X1  g793(.A(G227), .B1(new_n670), .B2(G14), .ZN(new_n1220));
  AND4_X1   g794(.A1(new_n900), .A2(new_n977), .A3(new_n1219), .A4(new_n1220), .ZN(G308));
  NAND4_X1  g795(.A1(new_n900), .A2(new_n977), .A3(new_n1219), .A4(new_n1220), .ZN(G225));
endmodule


