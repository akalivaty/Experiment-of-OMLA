//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT70), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n196));
  XOR2_X1   g010(.A(new_n196), .B(KEYINPUT22), .Z(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G119), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(KEYINPUT74), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT74), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(KEYINPUT23), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT75), .B(G110), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n203), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n202), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT76), .A3(new_n213), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(G125), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n221), .A2(KEYINPUT16), .A3(G140), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(G146), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n203), .A2(new_n207), .ZN(new_n229));
  INV_X1    g043(.A(G110), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n220), .A2(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n224), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n223), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n211), .A2(new_n212), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n236), .A3(KEYINPUT77), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT77), .B1(new_n228), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n199), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n199), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n188), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n243), .B2(KEYINPUT25), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(KEYINPUT25), .B2(new_n243), .ZN(new_n245));
  INV_X1    g059(.A(new_n239), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n237), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n238), .A2(new_n199), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n190), .A2(new_n188), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(KEYINPUT79), .A3(new_n251), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G119), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n204), .B2(G116), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(KEYINPUT69), .A3(G119), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT2), .B(G113), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n198), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G137), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT11), .A2(G134), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G137), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(G137), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(KEYINPUT11), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT11), .B1(new_n198), .B2(G134), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n198), .A2(G134), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n274), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n290));
  OAI22_X1  g104(.A1(new_n289), .A2(new_n290), .B1(KEYINPUT0), .B2(G128), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT65), .A2(G143), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT65), .A2(G143), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n224), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n224), .A2(G143), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n224), .A2(G143), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n293), .A2(new_n294), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(G146), .ZN(new_n302));
  INV_X1    g116(.A(new_n287), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n292), .A2(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n286), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT65), .B(G143), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n296), .B1(new_n306), .B2(new_n224), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n200), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT68), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n308), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n309), .A2(new_n312), .B1(new_n302), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(G134), .B1(new_n270), .B2(new_n272), .ZN(new_n315));
  OAI21_X1  g129(.A(G131), .B1(new_n315), .B2(new_n278), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n285), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n305), .B(KEYINPUT30), .C1(new_n314), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n283), .A2(new_n284), .A3(new_n274), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n284), .B1(new_n283), .B2(new_n274), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n299), .B1(new_n306), .B2(new_n224), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n323), .A2(new_n287), .B1(new_n307), .B2(new_n291), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n319), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n286), .A2(new_n304), .A3(KEYINPUT67), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n299), .B(new_n313), .C1(new_n306), .C2(new_n224), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n307), .A2(KEYINPUT68), .A3(new_n308), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n311), .B1(new_n298), .B2(new_n310), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n317), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n325), .A2(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n269), .B(new_n318), .C1(new_n332), .C2(KEYINPUT30), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n268), .A3(new_n305), .ZN(new_n335));
  INV_X1    g149(.A(G237), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n192), .A2(new_n194), .A3(G210), .A4(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n337), .B(KEYINPUT27), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT26), .ZN(new_n347));
  AOI21_X1  g161(.A(G101), .B1(new_n347), .B2(new_n341), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n333), .A2(new_n335), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT31), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n335), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n334), .A2(KEYINPUT28), .A3(new_n268), .A4(new_n305), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n332), .A2(new_n268), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n347), .A2(G101), .A3(new_n341), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT71), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n355), .A2(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n333), .A2(new_n349), .A3(new_n362), .A4(new_n335), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n351), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G472), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n257), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g182(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n364), .A2(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n333), .A2(new_n335), .ZN(new_n372));
  INV_X1    g186(.A(new_n349), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n359), .A2(new_n360), .ZN(new_n375));
  INV_X1    g189(.A(new_n356), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n353), .A4(new_n354), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n345), .A2(new_n348), .A3(new_n378), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n334), .A2(new_n305), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n269), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n353), .A2(new_n380), .A3(new_n382), .A4(new_n354), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT73), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n188), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n188), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n371), .A2(KEYINPUT32), .B1(new_n388), .B2(G472), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n256), .B1(new_n370), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G214), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G104), .ZN(new_n397));
  OR2_X1    g211(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n401), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT81), .B(G101), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n399), .ZN(new_n406));
  INV_X1    g220(.A(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n396), .A2(G104), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n397), .B2(new_n398), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n410), .A3(new_n343), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n268), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n259), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(G113), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G101), .B1(new_n407), .B2(new_n409), .ZN(new_n421));
  AND4_X1   g235(.A1(new_n265), .A2(new_n420), .A3(new_n411), .A4(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n395), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n415), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n414), .B1(new_n405), .B2(new_n411), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n269), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n411), .A2(new_n421), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n265), .A3(new_n420), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(new_n394), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n221), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n324), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n191), .A2(G224), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT88), .Z(new_n436));
  XNOR2_X1  g250(.A(new_n434), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n395), .C1(new_n416), .C2(new_n422), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(new_n188), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n394), .B(KEYINPUT8), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n420), .A2(new_n265), .B1(new_n411), .B2(new_n421), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n422), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n435), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(KEYINPUT89), .B2(new_n446), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n434), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n432), .A2(KEYINPUT7), .A3(new_n433), .A4(new_n435), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n445), .A2(new_n451), .A3(new_n455), .A4(new_n452), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n456), .A3(new_n430), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n441), .A2(new_n442), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n188), .A3(new_n440), .ZN(new_n459));
  INV_X1    g273(.A(new_n442), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n393), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n195), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(G902), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(G898), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n464), .A2(G952), .A3(new_n191), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT15), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G478), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n187), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n301), .A2(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n200), .A2(G143), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n276), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT97), .B1(new_n479), .B2(G116), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n258), .A3(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n258), .B2(G122), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(G107), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(G107), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT13), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n477), .B1(new_n476), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n306), .A2(new_n200), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT98), .B1(new_n490), .B2(KEYINPUT13), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n476), .A2(new_n492), .A3(new_n488), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n487), .B1(new_n495), .B2(G134), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n476), .A2(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G134), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n478), .ZN(new_n499));
  INV_X1    g313(.A(new_n486), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n483), .A2(KEYINPUT14), .B1(new_n258), .B2(G122), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n502));
  OAI21_X1  g316(.A(G107), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n475), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n494), .A2(new_n276), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n504), .B(new_n474), .C1(new_n507), .C2(new_n487), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT99), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n511), .B(G902), .C1(new_n506), .C2(new_n508), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n472), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n512), .A2(new_n472), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n192), .A2(new_n194), .A3(G214), .A4(new_n336), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n301), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n520), .A3(new_n301), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n195), .A2(G143), .A3(G214), .A4(new_n336), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n519), .A2(new_n522), .A3(new_n524), .A4(new_n521), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n219), .B(new_n224), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT94), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(new_n401), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(G131), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n519), .A2(new_n522), .A3(new_n284), .A4(new_n521), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n233), .A2(new_n223), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n533), .B2(new_n534), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n529), .B(new_n532), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n532), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n219), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n219), .A2(new_n542), .A3(KEYINPUT93), .ZN(new_n546));
  INV_X1    g360(.A(new_n219), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT19), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n545), .A2(new_n224), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n223), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n533), .B2(new_n535), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n540), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G475), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n188), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n539), .A2(new_n558), .A3(new_n552), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n539), .B2(new_n552), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n559), .A2(new_n560), .A3(new_n555), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n529), .B1(new_n536), .B2(new_n538), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n540), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n565), .B2(new_n539), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT96), .B(G475), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n516), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n470), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n330), .A2(new_n428), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n200), .B1(new_n295), .B2(KEYINPUT1), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT83), .B1(new_n573), .B2(new_n302), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT83), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT1), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n306), .B2(new_n224), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n323), .C1(new_n577), .C2(new_n200), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT82), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n327), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n302), .A2(KEYINPUT82), .A3(new_n313), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n574), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n428), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(KEYINPUT84), .A3(new_n428), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n572), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT12), .B1(new_n587), .B2(new_n322), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n582), .A2(KEYINPUT84), .A3(new_n428), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT84), .B1(new_n582), .B2(new_n428), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n589), .A2(new_n590), .B1(new_n330), .B2(new_n428), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT12), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n286), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n589), .B2(new_n590), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n413), .A2(new_n415), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n427), .A2(new_n594), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n596), .A2(new_n304), .B1(new_n330), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n322), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT85), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n588), .A2(new_n602), .A3(new_n593), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n195), .A2(G227), .ZN(new_n605));
  XOR2_X1   g419(.A(G110), .B(G140), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n322), .A2(KEYINPUT86), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT10), .B1(new_n585), .B2(new_n586), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n596), .A2(new_n304), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n330), .A2(new_n597), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n609), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n609), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n595), .A2(new_n598), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n607), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n608), .A2(G469), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n607), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n588), .A2(new_n621), .A3(new_n593), .A4(new_n599), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(KEYINPUT87), .B1(new_n617), .B2(new_n607), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n585), .A2(new_n586), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n613), .B1(new_n624), .B2(new_n594), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n591), .A2(new_n286), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n322), .A2(new_n625), .B1(new_n626), .B2(KEYINPUT12), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT87), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n621), .A4(new_n593), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G469), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n188), .ZN(new_n632));
  NAND2_X1  g446(.A1(G469), .A2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n620), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n571), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n391), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n343), .ZN(G3));
  AND2_X1   g452(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n364), .A2(new_n188), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n366), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n256), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n506), .A2(new_n508), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n506), .A2(KEYINPUT33), .A3(new_n508), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(G478), .A3(new_n188), .A4(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n509), .A2(G478), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n553), .A2(KEYINPUT95), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n539), .A2(new_n558), .A3(new_n552), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n554), .A3(new_n188), .A4(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(KEYINPUT20), .B1(new_n553), .B2(new_n556), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n652), .B1(new_n656), .B2(new_n568), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n470), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n645), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NAND2_X1  g475(.A1(new_n515), .A2(new_n569), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n458), .A2(new_n461), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n469), .B(KEYINPUT103), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n392), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n561), .B2(new_n562), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n655), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n559), .A2(new_n560), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n556), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n667), .A2(new_n668), .A3(new_n673), .A4(new_n670), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n662), .B(new_n665), .C1(new_n672), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n645), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n228), .A2(new_n236), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n251), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n245), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n366), .A3(new_n641), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n571), .A2(new_n634), .A3(new_n684), .A4(new_n635), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT37), .B(G110), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT104), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n366), .A2(new_n367), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT72), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n366), .A2(new_n257), .A3(new_n367), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n389), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n683), .A2(new_n462), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n692), .A2(new_n634), .A3(new_n635), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n468), .B1(new_n465), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n662), .B(new_n696), .C1(new_n672), .C2(new_n674), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n696), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n639), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n663), .B(KEYINPUT105), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT38), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n515), .B1(new_n656), .B2(new_n568), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n683), .A3(new_n393), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n375), .B1(new_n335), .B2(new_n382), .ZN(new_n708));
  INV_X1    g522(.A(new_n350), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n188), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n371), .A2(KEYINPUT32), .B1(G472), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n370), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT106), .Z(new_n713));
  NOR2_X1   g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n702), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT107), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n306), .ZN(G45));
  INV_X1    g531(.A(new_n696), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n652), .B(new_n718), .C1(new_n656), .C2(new_n568), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n693), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n639), .A2(new_n692), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  AOI21_X1  g537(.A(new_n631), .B1(new_n630), .B2(new_n188), .ZN(new_n724));
  AOI211_X1 g538(.A(G469), .B(G902), .C1(new_n623), .C2(new_n629), .ZN(new_n725));
  INV_X1    g539(.A(new_n635), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n390), .A3(new_n658), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND3_X1  g544(.A1(new_n675), .A2(new_n390), .A3(new_n727), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  INV_X1    g546(.A(new_n570), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n692), .A2(new_n469), .A3(new_n733), .A4(new_n683), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n630), .A2(new_n188), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n635), .A3(new_n632), .A4(new_n462), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n442), .B1(new_n441), .B2(new_n457), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n459), .A2(new_n460), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n392), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n740), .B1(new_n705), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n563), .A2(new_n569), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n462), .A2(new_n745), .A3(KEYINPUT108), .A4(new_n515), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n355), .B1(new_n269), .B2(new_n381), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n351), .B(new_n363), .C1(new_n748), .C2(new_n375), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n365), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n641), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n256), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n747), .A2(new_n727), .A3(new_n664), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  INV_X1    g569(.A(new_n751), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n720), .A2(new_n756), .A3(new_n683), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n755), .B1(new_n737), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n683), .A2(new_n641), .A3(new_n750), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n719), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n727), .A2(new_n760), .A3(KEYINPUT109), .A4(new_n462), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NAND3_X1  g577(.A1(new_n458), .A2(new_n461), .A3(new_n392), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n256), .B(new_n764), .C1(new_n370), .C2(new_n389), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n608), .A2(KEYINPUT111), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n621), .B1(new_n601), .B2(new_n603), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n618), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n769), .A3(G469), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n633), .B(KEYINPUT110), .Z(new_n771));
  AOI21_X1  g585(.A(G902), .B1(new_n623), .B2(new_n629), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n631), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n726), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n774), .A3(new_n720), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n256), .B1(new_n389), .B2(new_n689), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n719), .A2(new_n776), .A3(new_n764), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND2_X1  g596(.A1(new_n672), .A2(new_n674), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  INV_X1    g598(.A(new_n662), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n718), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n765), .A2(new_n786), .A3(new_n774), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n697), .A2(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND3_X1  g604(.A1(new_n766), .A2(new_n769), .A3(KEYINPUT45), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n767), .A2(new_n618), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n791), .B(G469), .C1(KEYINPUT45), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n771), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n632), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n745), .B1(new_n651), .B2(new_n650), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n799), .B2(KEYINPUT113), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n642), .A3(new_n683), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n806), .A3(new_n764), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n798), .A2(new_n807), .A3(new_n635), .A4(new_n700), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  OAI21_X1  g623(.A(new_n635), .B1(new_n796), .B2(new_n797), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n635), .C1(new_n796), .C2(new_n797), .ZN(new_n813));
  INV_X1    g627(.A(new_n256), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n692), .A2(new_n814), .A3(new_n719), .A4(new_n764), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  AND3_X1   g632(.A1(new_n801), .A2(new_n468), .A3(new_n802), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n752), .ZN(new_n820));
  OAI211_X1 g634(.A(G952), .B(new_n191), .C1(new_n820), .C2(new_n737), .ZN(new_n821));
  INV_X1    g635(.A(new_n764), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n727), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n814), .A2(new_n825), .A3(new_n468), .A4(new_n713), .ZN(new_n826));
  INV_X1    g640(.A(new_n657), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n825), .A2(new_n819), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT48), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n829), .A2(new_n830), .A3(new_n778), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n829), .B2(new_n778), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n759), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n704), .A2(new_n392), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n727), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n839), .A2(new_n820), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n839), .B2(new_n820), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n745), .A2(new_n652), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n841), .A2(new_n842), .B1(new_n826), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n837), .A2(KEYINPUT51), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n811), .A2(new_n813), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n724), .A2(new_n725), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n635), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n820), .A2(new_n764), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n833), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n822), .A2(new_n683), .A3(new_n718), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n770), .A2(new_n773), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n751), .A2(new_n657), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n635), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n516), .A2(new_n569), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n672), .B2(new_n674), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n692), .A3(new_n635), .A4(new_n634), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n854), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n563), .A2(new_n515), .A3(new_n569), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n665), .B1(new_n862), .B2(new_n657), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n634), .A3(new_n635), .A4(new_n643), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n685), .C1(new_n391), .C2(new_n636), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n781), .A3(new_n789), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n783), .A2(new_n462), .A3(new_n785), .A4(new_n664), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n847), .A2(new_n692), .A3(new_n814), .A4(new_n635), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n728), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n847), .A2(new_n635), .A3(new_n664), .A4(new_n752), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n744), .A2(new_n746), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(new_n734), .B2(new_n737), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n868), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n390), .B(new_n727), .C1(new_n675), .C2(new_n658), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n738), .A3(KEYINPUT115), .A4(new_n753), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n683), .A2(new_n696), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n774), .A2(new_n712), .A3(new_n747), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n762), .A2(new_n698), .A3(new_n722), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n758), .A2(new_n761), .B1(new_n694), .B2(new_n697), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n722), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n853), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n882), .A2(new_n890), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n777), .A2(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n875), .A3(new_n877), .A4(new_n866), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT53), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n884), .A2(new_n886), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n853), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(new_n867), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n871), .A2(new_n874), .A3(new_n853), .ZN(new_n904));
  INV_X1    g718(.A(new_n893), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n891), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n852), .A2(new_n899), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n837), .A2(new_n844), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n851), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n849), .A2(KEYINPUT118), .A3(new_n850), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT51), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n908), .A2(new_n913), .B1(G952), .B2(G953), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n799), .A2(new_n814), .A3(new_n635), .A4(new_n392), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n704), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n847), .B(KEYINPUT49), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n713), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n195), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n879), .B2(new_n887), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n895), .A2(new_n904), .A3(new_n866), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n892), .B2(new_n893), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n188), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n431), .A2(new_n439), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n437), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT121), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT55), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n921), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n927), .B2(new_n932), .ZN(G51));
  NOR3_X1   g748(.A1(new_n925), .A2(new_n188), .A3(new_n793), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT54), .B1(new_n922), .B2(new_n924), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(KEYINPUT122), .A3(new_n907), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(KEYINPUT54), .C1(new_n922), .C2(new_n924), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n771), .B(KEYINPUT57), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n630), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n935), .B1(new_n942), .B2(KEYINPUT123), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n944), .A3(new_n630), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n920), .B1(new_n943), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n669), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n920), .ZN(G60));
  AND2_X1   g765(.A1(new_n648), .A2(new_n649), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n899), .A2(new_n907), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n952), .A2(new_n937), .A3(new_n939), .A4(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n920), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n925), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(new_n249), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n681), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n921), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n921), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G66));
  INV_X1    g782(.A(G224), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n466), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n878), .A2(new_n865), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n195), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n928), .B1(G898), .B2(new_n195), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  OAI21_X1  g790(.A(new_n318), .B1(new_n332), .B2(KEYINPUT30), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n195), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n885), .A2(new_n722), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n715), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n715), .A2(new_n985), .A3(new_n982), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n657), .A2(new_n862), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n639), .A2(new_n765), .A3(new_n700), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n817), .A2(new_n808), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n981), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n980), .B1(new_n695), .B2(new_n463), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n747), .A2(new_n778), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n798), .A2(new_n635), .A3(new_n700), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n982), .A2(new_n895), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n817), .A2(new_n808), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n995), .B1(new_n999), .B2(new_n195), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT126), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n195), .B(new_n980), .C1(new_n989), .C2(new_n991), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n999), .A2(new_n195), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n995), .ZN(new_n1005));
  INV_X1    g819(.A(G227), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n463), .B1(new_n1006), .B2(new_n695), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1001), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  OR2_X1    g824(.A1(new_n999), .A2(new_n972), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  AOI211_X1 g827(.A(new_n349), .B(new_n372), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n372), .A2(new_n349), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n989), .A2(new_n991), .A3(new_n972), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1016), .B2(new_n1013), .ZN(new_n1017));
  INV_X1    g831(.A(new_n374), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1013), .B1(new_n1018), .B2(new_n709), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT127), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n898), .A2(new_n1020), .ZN(new_n1021));
  NOR4_X1   g835(.A1(new_n1014), .A2(new_n1017), .A3(new_n920), .A4(new_n1021), .ZN(G57));
endmodule


