//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(new_n195), .C1(new_n196), .C2(KEYINPUT23), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT75), .B(G110), .Z(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n200));
  OAI22_X1  g014(.A1(new_n197), .A2(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT16), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n205), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n201), .B(new_n208), .C1(G146), .C2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n197), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n211));
  INV_X1    g025(.A(new_n208), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n206), .B2(new_n207), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT76), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n215), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n188), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n191), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT25), .B(new_n188), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n190), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n223), .A2(G902), .A3(new_n189), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(G472), .A2(G902), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT0), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(new_n192), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G143), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n237), .A2(KEYINPUT64), .A3(G146), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT64), .B1(new_n237), .B2(G146), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n234), .B(new_n236), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n192), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT65), .A2(G131), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT65), .A2(G131), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(new_n251), .A3(new_n249), .A4(new_n252), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n254), .A2(new_n258), .A3(KEYINPUT70), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n254), .B2(new_n258), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n246), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G128), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n236), .B(new_n264), .C1(new_n238), .C2(new_n239), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(G143), .B2(new_n235), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n243), .B1(new_n266), .B2(new_n192), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G134), .B(G137), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT66), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n248), .A2(G137), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n250), .A2(G134), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n272), .B(G131), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n258), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n277), .A3(KEYINPUT30), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n265), .A2(new_n267), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n258), .A2(new_n271), .A3(new_n283), .A4(new_n275), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n254), .A2(new_n258), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n246), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT2), .B(G113), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G116), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G119), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT69), .B(G116), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(G119), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n292), .B1(new_n296), .B2(KEYINPUT68), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(G119), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n293), .B2(G119), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n291), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n261), .A2(new_n277), .A3(KEYINPUT71), .A4(KEYINPUT30), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n280), .A2(new_n290), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT27), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G101), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n305), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n261), .A2(new_n313), .A3(new_n277), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n307), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT31), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n307), .A2(KEYINPUT31), .A3(new_n312), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n314), .A2(new_n320), .B1(new_n288), .B2(new_n305), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n261), .A2(new_n313), .A3(new_n277), .A4(KEYINPUT28), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n312), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n232), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n320), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  INV_X1    g142(.A(new_n314), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n313), .B1(new_n261), .B2(new_n277), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n288), .A2(new_n305), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n327), .A2(new_n336), .A3(new_n312), .A4(new_n322), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n321), .A2(new_n339), .A3(new_n312), .A4(new_n322), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(new_n333), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n312), .B1(new_n307), .B2(new_n314), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n335), .B(new_n188), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n326), .A2(KEYINPUT32), .B1(G472), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n317), .A2(new_n318), .B1(new_n324), .B2(new_n323), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n232), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n230), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT9), .B(G234), .ZN(new_n349));
  OAI21_X1  g163(.A(G221), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n259), .A2(new_n260), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n361), .A3(G104), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n358), .B(new_n366), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n369), .A3(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n246), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT78), .B(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n357), .B1(new_n372), .B2(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n282), .A2(new_n374), .A3(KEYINPUT10), .A4(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n378), .B(KEYINPUT1), .C1(new_n237), .C2(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G128), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n237), .A2(G146), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT64), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n242), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n237), .A2(KEYINPUT64), .A3(G146), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n377), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(KEYINPUT80), .C1(new_n381), .C2(new_n380), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n265), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n374), .A2(new_n367), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT10), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n353), .B1(new_n376), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n353), .C1(new_n376), .C2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G140), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n216), .A2(G227), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n374), .A2(new_n367), .ZN(new_n403));
  INV_X1    g217(.A(new_n265), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n389), .B1(new_n381), .B2(new_n380), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n377), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n406), .B2(new_n390), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n371), .B(new_n375), .C1(new_n407), .C2(KEYINPUT10), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n402), .B1(new_n408), .B2(new_n353), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n376), .A2(new_n393), .A3(new_n353), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT12), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n254), .B2(new_n258), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n403), .A2(new_n268), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n391), .A2(new_n392), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n352), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n418), .B2(KEYINPUT12), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n398), .A2(new_n410), .B1(new_n420), .B2(new_n401), .ZN(new_n421));
  OAI21_X1  g235(.A(G469), .B1(new_n421), .B2(G902), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n408), .A2(new_n353), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n395), .B2(new_n397), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n353), .B1(new_n407), .B2(new_n415), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n414), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n425), .A2(new_n412), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n424), .A2(new_n402), .B1(new_n409), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n188), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n351), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n368), .A2(new_n305), .A3(new_n370), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n296), .A2(new_n292), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n294), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(G113), .B(new_n435), .C1(new_n302), .C2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n392), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT82), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n240), .A2(new_n245), .A3(G125), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(G125), .B1(new_n265), .B2(new_n267), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n282), .A2(new_n204), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT83), .B1(new_n452), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT84), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n216), .A2(G224), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(KEYINPUT83), .A3(new_n447), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n454), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(new_n454), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n444), .B(new_n446), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n452), .B(new_n447), .C1(KEYINPUT85), .C2(new_n456), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n436), .A2(new_n433), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n403), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n437), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n440), .B(KEYINPUT8), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n466), .A2(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n472), .B2(new_n443), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n474), .B(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G214), .B1(G237), .B2(G902), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G478), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n298), .A2(new_n300), .A3(G122), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n293), .A2(G122), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G107), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT95), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n484), .A2(new_n486), .ZN(new_n490));
  XOR2_X1   g304(.A(G128), .B(G143), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G134), .ZN(new_n492));
  XNOR2_X1  g306(.A(G128), .B(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n248), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n490), .A2(new_n372), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n295), .A2(KEYINPUT14), .A3(G122), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n497), .A3(G107), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n237), .A3(G128), .ZN(new_n502));
  OAI211_X1 g316(.A(G134), .B(new_n502), .C1(new_n491), .C2(new_n501), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n490), .A2(new_n372), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n484), .A2(new_n372), .A3(new_n486), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n503), .B(new_n494), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n349), .A2(new_n187), .A3(G953), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n506), .A3(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n483), .B1(new_n512), .B2(new_n188), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n500), .A2(new_n506), .A3(new_n508), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n508), .B1(new_n500), .B2(new_n506), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n483), .B(new_n188), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n482), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n481), .A3(G478), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G902), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n209), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT89), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(G146), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n203), .A2(new_n205), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n235), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n523), .A2(new_n526), .A3(G146), .A4(new_n524), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n270), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n308), .A2(G214), .B1(new_n533), .B2(G143), .ZN(new_n534));
  INV_X1    g348(.A(G214), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n535), .A2(G237), .A3(G953), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n237), .A2(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n534), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n532), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n533), .A2(G143), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n237), .A2(KEYINPUT88), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n536), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G237), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n216), .A3(G214), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n538), .ZN(new_n548));
  AND4_X1   g362(.A1(new_n541), .A2(new_n545), .A3(new_n532), .A4(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n529), .B(new_n530), .C1(new_n542), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n257), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n547), .B1(new_n537), .B2(new_n538), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(new_n534), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n257), .A3(new_n548), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n212), .A2(new_n213), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n545), .A2(new_n548), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT17), .A3(new_n551), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(G113), .B(G122), .Z(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G104), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n550), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n550), .B2(new_n560), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n521), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n550), .A2(new_n560), .A3(new_n562), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n529), .A2(new_n530), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n558), .A2(KEYINPUT91), .B1(new_n531), .B2(new_n270), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n540), .A2(new_n541), .A3(new_n532), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n523), .A2(KEYINPUT19), .A3(new_n524), .ZN(new_n572));
  OR2_X1    g386(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n573));
  NAND2_X1  g387(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n527), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n235), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n212), .B1(new_n553), .B2(new_n555), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n568), .A2(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n567), .B1(new_n578), .B2(new_n562), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT20), .ZN(new_n581));
  NOR2_X1   g395(.A1(G475), .A2(G902), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT93), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(new_n576), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n562), .B1(new_n550), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n581), .B(new_n584), .C1(new_n563), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n579), .B2(new_n584), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n566), .B(new_n585), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G952), .ZN(new_n593));
  AOI211_X1 g407(.A(G953), .B(new_n593), .C1(G234), .C2(G237), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n216), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n520), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n479), .A2(new_n480), .A3(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n348), .A2(new_n431), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n366), .ZN(G3));
  NAND2_X1  g415(.A1(new_n319), .A2(new_n325), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n188), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n326), .B1(new_n603), .B2(G472), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n229), .A3(new_n431), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n474), .A2(new_n475), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n463), .A2(new_n473), .A3(new_n476), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n480), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n592), .ZN(new_n609));
  INV_X1    g423(.A(G478), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n224), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT33), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n510), .B2(new_n511), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n188), .B1(new_n514), .B2(new_n515), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n610), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR4_X1   g434(.A1(new_n605), .A2(new_n597), .A3(new_n608), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n520), .A2(new_n566), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n590), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n563), .A2(new_n587), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(new_n583), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n579), .A2(new_n584), .A3(new_n590), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n597), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n579), .A2(KEYINPUT97), .A3(new_n584), .A4(new_n590), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n625), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n605), .A2(new_n608), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT35), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n215), .B(new_n640), .Z(new_n641));
  NOR2_X1   g455(.A1(new_n189), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n227), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  INV_X1    g460(.A(new_n227), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n643), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n599), .A2(new_n604), .A3(new_n431), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  NAND3_X1  g467(.A1(new_n602), .A2(KEYINPUT32), .A3(new_n231), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n343), .A2(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n347), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n594), .B1(new_n595), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n565), .B2(G475), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n520), .A2(new_n633), .A3(new_n631), .A4(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n658), .B1(new_n608), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n631), .A2(new_n633), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n616), .A2(KEYINPUT96), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n665), .A2(new_n516), .B1(new_n481), .B2(G478), .ZN(new_n666));
  INV_X1    g480(.A(new_n519), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n476), .B1(new_n463), .B2(new_n473), .ZN(new_n670));
  INV_X1    g484(.A(new_n480), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(KEYINPUT99), .A3(new_n607), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n663), .A2(new_n673), .A3(new_n431), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n657), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n192), .ZN(G30));
  XOR2_X1   g490(.A(new_n660), .B(KEYINPUT39), .Z(new_n677));
  AND2_X1   g491(.A1(new_n431), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  INV_X1    g493(.A(G472), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n315), .B2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n654), .B(new_n347), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n479), .B(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n520), .A2(new_n592), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n650), .A2(new_n671), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n679), .A2(new_n683), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n463), .A2(new_n473), .A3(new_n476), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n690), .A2(new_n670), .A3(new_n671), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n615), .A2(new_n617), .ZN(new_n692));
  INV_X1    g506(.A(new_n660), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n592), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT100), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n592), .A2(new_n692), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n695), .A3(KEYINPUT101), .A4(new_n697), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n431), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n689), .B1(new_n702), .B2(new_n657), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n422), .A2(new_n430), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n350), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n699), .B2(new_n698), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n344), .A2(new_n347), .B1(new_n646), .B2(new_n649), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(KEYINPUT102), .A3(new_n707), .A4(new_n701), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND4_X1  g524(.A1(new_n656), .A2(new_n229), .A3(new_n632), .A4(new_n619), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n409), .A2(new_n427), .ZN(new_n712));
  INV_X1    g526(.A(new_n397), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n396), .B1(new_n408), .B2(new_n353), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n411), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n712), .B1(new_n715), .B2(new_n401), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(new_n224), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT103), .A3(new_n430), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n719), .B(G469), .C1(new_n716), .C2(new_n224), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n350), .A3(new_n691), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  AOI211_X1 g539(.A(new_n351), .B(new_n608), .C1(new_n718), .C2(new_n720), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n348), .A4(new_n635), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n656), .A2(new_n635), .A3(new_n229), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT104), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  NAND3_X1  g546(.A1(new_n656), .A2(new_n598), .A3(new_n650), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n194), .ZN(G21));
  NAND3_X1  g549(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n324), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n232), .B1(new_n319), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n603), .B2(G472), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n685), .A2(new_n597), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n229), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n722), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(G122), .Z(G24));
  AND2_X1   g557(.A1(new_n695), .A2(new_n697), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n739), .A2(new_n744), .A3(new_n650), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n722), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n204), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n716), .A2(G469), .A3(new_n224), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n398), .A2(new_n410), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n420), .A2(new_n401), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n429), .B1(new_n752), .B2(new_n521), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n748), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n479), .A2(new_n671), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n422), .A2(new_n430), .A3(KEYINPUT105), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n350), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n656), .A2(new_n229), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n695), .A2(new_n697), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n350), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n347), .A2(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n347), .A2(KEYINPUT106), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n344), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n229), .A3(new_n765), .A4(new_n744), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n761), .B1(new_n766), .B2(KEYINPUT42), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT107), .B(G131), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G33));
  AND3_X1   g583(.A1(new_n422), .A2(new_n430), .A3(KEYINPUT105), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT105), .B1(new_n422), .B2(new_n430), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n771), .A3(new_n351), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n662), .B(KEYINPUT108), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n348), .A3(new_n755), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n348), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(new_n755), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n618), .A2(new_n592), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(KEYINPUT110), .B2(KEYINPUT43), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n618), .B2(new_n592), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n650), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(new_n604), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n421), .A2(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n421), .A2(KEYINPUT45), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(G469), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(G469), .A2(G902), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT46), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n749), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(KEYINPUT46), .A3(new_n794), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n351), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n677), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  OR2_X1    g615(.A1(new_n795), .A2(new_n749), .ZN(new_n802));
  INV_X1    g616(.A(new_n797), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n350), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n780), .A2(new_n656), .A3(new_n229), .A4(new_n759), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT111), .B(G140), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G42));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n813));
  NOR2_X1   g627(.A1(G952), .A2(G953), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n757), .A2(new_n745), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n780), .A2(new_n705), .A3(new_n520), .A4(new_n664), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n707), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n767), .A2(new_n778), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n645), .A2(new_n660), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n772), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n754), .A2(new_n350), .A3(new_n756), .A4(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n608), .A2(new_n685), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n823), .A3(new_n683), .A4(new_n824), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n722), .A2(new_n745), .B1(new_n657), .B2(new_n674), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n709), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n703), .B2(new_n708), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n825), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n818), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n479), .A2(new_n480), .A3(new_n632), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n620), .A2(KEYINPUT115), .B1(new_n836), .B2(new_n624), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n479), .A2(new_n480), .A3(new_n632), .A4(new_n619), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n835), .A2(new_n837), .B1(KEYINPUT115), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n651), .B1(new_n839), .B2(new_n605), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n600), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n722), .B1(new_n711), .B2(new_n741), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n734), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n731), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n731), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n833), .B2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n767), .A2(new_n778), .A3(new_n817), .ZN(new_n851));
  AND4_X1   g665(.A1(KEYINPUT52), .A2(new_n709), .A3(new_n827), .A4(new_n825), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(new_n831), .B2(new_n825), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n841), .A2(KEYINPUT53), .A3(new_n731), .A4(new_n844), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n850), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n731), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT114), .B1(new_n844), .B2(new_n731), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n841), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n859), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n833), .A2(new_n849), .A3(KEYINPUT53), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n739), .A2(new_n229), .ZN(new_n867));
  INV_X1    g681(.A(new_n594), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n782), .B2(new_n784), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n780), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n721), .A2(new_n351), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n806), .A2(new_n807), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n721), .A2(new_n350), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n780), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n683), .A2(new_n230), .A3(new_n868), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n609), .A3(new_n878), .A4(new_n618), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n650), .A3(new_n739), .A4(new_n869), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  INV_X1    g698(.A(new_n870), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n876), .A2(new_n684), .A3(new_n480), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT50), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT50), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n881), .A2(new_n882), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n875), .A2(new_n883), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n229), .A2(new_n877), .A3(new_n765), .A4(new_n869), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(KEYINPUT48), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(KEYINPUT48), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n877), .A2(new_n619), .A3(new_n878), .ZN(new_n897));
  OAI211_X1 g711(.A(G952), .B(new_n216), .C1(new_n870), .C2(new_n722), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n889), .A2(new_n890), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n881), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(KEYINPUT119), .A3(new_n881), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT118), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT118), .B1(new_n872), .B2(new_n874), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n884), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n814), .B1(new_n866), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n721), .B(KEYINPUT49), .Z(new_n911));
  NAND4_X1  g725(.A1(new_n781), .A2(new_n229), .A3(new_n350), .A4(new_n480), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT112), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n683), .A2(new_n911), .A3(new_n684), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT113), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n813), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n915), .ZN(new_n917));
  INV_X1    g731(.A(new_n864), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n918), .B2(new_n850), .ZN(new_n919));
  INV_X1    g733(.A(new_n855), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n833), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n863), .A2(new_n858), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n909), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT121), .B(new_n917), .C1(new_n923), .C2(new_n814), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n924), .ZN(G75));
  NAND2_X1  g739(.A1(new_n863), .A2(new_n921), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n224), .A3(new_n476), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n444), .A2(new_n446), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n929), .A2(new_n461), .A3(new_n462), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n463), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n927), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n927), .B2(new_n928), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n216), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G51));
  XOR2_X1   g750(.A(new_n794), .B(KEYINPUT57), .Z(new_n937));
  AOI21_X1  g751(.A(new_n858), .B1(new_n863), .B2(new_n921), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n922), .B1(new_n938), .B2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n940), .B(new_n858), .C1(new_n863), .C2(new_n921), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n428), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n926), .A2(new_n224), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(new_n793), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n943), .B2(new_n945), .ZN(G54));
  NAND2_X1  g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n627), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n935), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n944), .A2(new_n627), .A3(new_n947), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G60));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  NOR2_X1   g768(.A1(new_n866), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n612), .A2(new_n614), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n939), .A2(new_n941), .ZN(new_n958));
  INV_X1    g772(.A(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n957), .A2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n926), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n223), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n926), .A2(new_n641), .A3(new_n964), .ZN(new_n967));
  NOR2_X1   g781(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n935), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G66));
  INV_X1    g786(.A(new_n596), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n216), .B1(new_n973), .B2(G224), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n862), .B2(new_n216), .ZN(new_n975));
  INV_X1    g789(.A(G898), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n929), .B1(new_n976), .B2(G953), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  AOI21_X1  g792(.A(KEYINPUT62), .B1(new_n687), .B2(new_n831), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n687), .A2(new_n831), .A3(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n620), .B1(new_n624), .B2(new_n836), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n348), .A2(new_n678), .A3(new_n755), .A4(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n982), .A2(new_n800), .A3(new_n810), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n216), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n280), .A2(new_n290), .A3(new_n306), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n572), .A2(new_n575), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n216), .B1(G227), .B2(G900), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n765), .A2(new_n229), .A3(new_n824), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n799), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n800), .A2(new_n810), .A3(new_n831), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n767), .A2(new_n778), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n994), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n991), .A2(new_n993), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(KEYINPUT125), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1004), .B(new_n994), .C1(new_n999), .C2(G953), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1003), .A2(new_n990), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1002), .B1(new_n1006), .B2(new_n993), .ZN(G72));
  XNOR2_X1  g821(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n680), .A2(new_n521), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n999), .B2(new_n862), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n307), .A2(new_n314), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT127), .Z(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n324), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1013), .A2(new_n324), .ZN(new_n1017));
  OAI221_X1 g831(.A(new_n1011), .B1(new_n1017), .B2(new_n342), .C1(new_n918), .C2(new_n850), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1011), .B1(new_n985), .B2(new_n862), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n312), .A3(new_n1014), .ZN(new_n1020));
  AND4_X1   g834(.A1(new_n949), .A2(new_n1016), .A3(new_n1018), .A4(new_n1020), .ZN(G57));
endmodule


