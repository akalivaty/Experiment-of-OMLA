//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n451), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT70), .B(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n461), .A3(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n473), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI211_X1 g054(.A(KEYINPUT71), .B(new_n469), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n465), .B1(new_n472), .B2(new_n480), .ZN(G160));
  INV_X1    g056(.A(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n462), .A2(KEYINPUT72), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n462), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n485), .B(new_n486), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G138), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n478), .A2(new_n495), .B1(KEYINPUT73), .B2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(new_n495), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n462), .A2(new_n497), .A3(new_n461), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n473), .A2(new_n475), .A3(G126), .ZN(new_n501));
  NAND2_X1  g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G2105), .B1(G102), .B2(new_n468), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G50), .ZN(new_n512));
  INV_X1    g087(.A(new_n509), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(G50), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT75), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(new_n518), .A3(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G88), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n517), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND2_X1  g104(.A1(new_n520), .A2(new_n522), .ZN(new_n530));
  INV_X1    g105(.A(new_n519), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n523), .A2(G89), .A3(new_n524), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT76), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(G51), .A2(new_n510), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n523), .A2(G89), .A3(new_n524), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n533), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(G168));
  XOR2_X1   g121(.A(KEYINPUT78), .B(G52), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n510), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n523), .A2(new_n524), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n523), .B2(G64), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI211_X1 g130(.A(KEYINPUT77), .B(new_n552), .C1(new_n523), .C2(G64), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n551), .B1(new_n557), .B2(G651), .ZN(G171));
  AOI22_X1  g133(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n527), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n510), .A2(G43), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n549), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  AOI22_X1  g145(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n527), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n510), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n523), .A2(new_n524), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G91), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(G299));
  OR2_X1    g152(.A1(new_n553), .A2(new_n554), .ZN(new_n578));
  INV_X1    g153(.A(new_n556), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(new_n579), .A3(G651), .ZN(new_n580));
  INV_X1    g155(.A(new_n551), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G301));
  AND3_X1   g157(.A1(new_n541), .A2(KEYINPUT79), .A3(new_n545), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT79), .B1(new_n541), .B2(new_n545), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n583), .A2(new_n584), .ZN(G286));
  OAI21_X1  g160(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n510), .A2(G49), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n549), .ZN(G288));
  AND2_X1   g164(.A1(new_n523), .A2(G61), .ZN(new_n590));
  AND2_X1   g165(.A1(G73), .A2(G543), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT80), .B(G651), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n510), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n549), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n591), .B1(new_n523), .B2(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n527), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n592), .A2(new_n596), .A3(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n527), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n575), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n575), .A2(new_n606), .A3(G92), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT10), .B1(new_n549), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n510), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n527), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n605), .B1(G868), .B2(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XNOR2_X1  g192(.A(G299), .B(KEYINPUT81), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(new_n564), .ZN(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n614), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(new_n624), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT82), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n462), .A2(new_n468), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n638), .B(new_n639), .C1(G111), .C2(new_n461), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n483), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n488), .A2(new_n489), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G135), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT84), .Z(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n634), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n683), .C2(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT85), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G26), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT92), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n643), .A2(G140), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT91), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n484), .A2(G128), .ZN(new_n700));
  OAI221_X1 g275(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n697), .B1(new_n703), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G2067), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n694), .A2(G33), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT25), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(new_n461), .ZN(new_n712));
  INV_X1    g287(.A(G139), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n712), .C1(new_n713), .C2(new_n490), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT93), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n707), .B1(new_n715), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2072), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(G164), .A2(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G27), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G11), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n694), .B1(new_n724), .B2(G28), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(G28), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n726), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n694), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G160), .B2(new_n694), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(G2084), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G2084), .B2(new_n735), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n718), .A2(new_n722), .A3(new_n723), .A4(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G5), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G171), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G168), .B2(G16), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G1966), .Z(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(G16), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n564), .B2(new_n748), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1341), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n743), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n739), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n614), .B2(new_n739), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1348), .ZN(new_n755));
  NOR4_X1   g330(.A1(new_n706), .A2(new_n738), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n716), .A2(new_n717), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n748), .A2(KEYINPUT23), .A3(G20), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n759));
  INV_X1    g334(.A(G20), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n747), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G299), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n758), .B(new_n761), .C1(new_n762), .C2(new_n739), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n720), .A2(new_n721), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n644), .A2(G29), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n756), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n739), .A2(G23), .ZN(new_n770));
  INV_X1    g345(.A(G288), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n739), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT33), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1976), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n748), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n748), .ZN(new_n776));
  INV_X1    g351(.A(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n739), .A2(G6), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G305), .B2(G16), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G1981), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(G1981), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT89), .B(KEYINPUT32), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n774), .A2(new_n778), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT90), .B1(new_n787), .B2(KEYINPUT34), .ZN(new_n789));
  MUX2_X1   g364(.A(G24), .B(G290), .S(new_n747), .Z(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1986), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n694), .A2(G25), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n643), .A2(G131), .B1(G119), .B2(new_n484), .ZN(new_n793));
  OAI221_X1 g368(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT86), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT87), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(new_n694), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n768), .B1(new_n769), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n769), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n694), .A2(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n694), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT29), .Z(new_n807));
  INV_X1    g382(.A(G2090), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n803), .A2(new_n804), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT26), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n643), .B2(G141), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n468), .A2(G105), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n484), .A2(G129), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G32), .B(new_n818), .S(G29), .Z(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT94), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT27), .B(G1996), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n812), .A2(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  OR2_X1    g399(.A1(new_n559), .A2(new_n527), .ZN(new_n825));
  INV_X1    g400(.A(new_n563), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n523), .A2(G67), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n527), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n510), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n549), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n825), .B(new_n826), .C1(new_n829), .C2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n829), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n834), .B(new_n835), .C1(new_n560), .C2(new_n563), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n614), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT97), .Z(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(KEYINPUT39), .C2(new_n840), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n834), .A2(new_n835), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(G145));
  XOR2_X1   g425(.A(new_n492), .B(KEYINPUT99), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G160), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n644), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n644), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n797), .ZN(new_n856));
  INV_X1    g431(.A(new_n797), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n818), .B(G164), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n703), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n715), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n643), .A2(G142), .B1(G130), .B2(new_n484), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n461), .A2(G118), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT100), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n632), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n862), .B(new_n869), .C1(new_n861), .C2(new_n714), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n861), .A2(new_n715), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n861), .A2(new_n714), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n859), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n856), .A3(new_n858), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g454(.A(G290), .B(G288), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  XNOR2_X1  g458(.A(G305), .B(G303), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n881), .A3(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n889), .B2(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n833), .A2(new_n836), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n627), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(KEYINPUT101), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n572), .A2(new_n574), .A3(new_n898), .A4(new_n576), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n626), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n762), .A2(new_n898), .A3(new_n614), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n907), .A3(new_n901), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n894), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n894), .A2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n847), .A2(new_n624), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(G331));
  XOR2_X1   g493(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  OAI21_X1  g495(.A(G171), .B1(new_n583), .B2(new_n584), .ZN(new_n921));
  NAND2_X1  g496(.A1(G301), .A2(G168), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(new_n895), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n895), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n895), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n903), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n909), .B(new_n910), .C1(new_n923), .C2(new_n924), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(KEYINPUT107), .A3(new_n903), .A4(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(new_n888), .ZN(new_n934));
  INV_X1    g509(.A(new_n888), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n930), .A2(new_n935), .A3(new_n931), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n877), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n925), .A2(new_n927), .B1(new_n908), .B2(new_n905), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n923), .A2(new_n924), .A3(new_n902), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n888), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n936), .A2(new_n941), .A3(new_n942), .A4(new_n877), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n919), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n936), .A2(new_n941), .A3(new_n877), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n933), .A2(new_n888), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(new_n942), .A3(new_n877), .A4(new_n936), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT44), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(new_n943), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n877), .A3(new_n936), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n951), .B(new_n952), .C1(new_n955), .C2(new_n919), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n505), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n463), .A2(new_n464), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n482), .ZN(new_n962));
  INV_X1    g537(.A(new_n480), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT71), .B1(new_n466), .B2(new_n469), .ZN(new_n964));
  OAI211_X1 g539(.A(G40), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n703), .A2(G2067), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n699), .A2(new_n705), .A3(new_n702), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n818), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n857), .A2(new_n799), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n797), .A2(new_n800), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(G290), .A2(G1986), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n966), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(G1384), .C1(new_n500), .C2(new_n504), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n959), .A2(new_n981), .A3(new_n965), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n721), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n505), .A2(new_n958), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n500), .B2(new_n504), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n965), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n742), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n983), .A2(new_n996), .A3(new_n984), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n986), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT124), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n984), .B1(new_n983), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n999), .B2(new_n983), .ZN(new_n1001));
  AOI21_X1  g576(.A(G301), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n982), .A2(KEYINPUT53), .A3(new_n721), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n986), .A2(new_n995), .A3(new_n997), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n979), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n998), .A2(G301), .A3(new_n1001), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n979), .B1(new_n1004), .B2(G171), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  INV_X1    g585(.A(G2084), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n988), .A2(new_n1011), .A3(new_n992), .A4(new_n993), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n982), .B2(G1966), .ZN(new_n1013));
  INV_X1    g588(.A(G168), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1012), .B(G168), .C1(new_n982), .C2(G1966), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1010), .B1(new_n1016), .B2(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT123), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(new_n1022), .C1(new_n1017), .C2(new_n1015), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT55), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n965), .B1(new_n1033), .B2(new_n989), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n987), .A2(new_n990), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n808), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n982), .B2(G1971), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1032), .B1(new_n1037), .B2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  AND3_X1   g614(.A1(G303), .A2(G8), .A3(new_n1030), .ZN(new_n1040));
  AOI22_X1  g615(.A1(G303), .A2(G8), .B1(new_n1026), .B2(KEYINPUT55), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1028), .A2(KEYINPUT111), .A3(new_n1031), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n982), .A2(G1971), .B1(new_n994), .B2(G2090), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n575), .A2(G87), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(G1976), .A3(new_n586), .A4(new_n587), .ZN(new_n1048));
  OAI211_X1 g623(.A(G8), .B(new_n1048), .C1(new_n987), .C2(new_n965), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n771), .A2(G1976), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1049), .A2(KEYINPUT52), .A3(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT113), .B(G1981), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n592), .A2(new_n596), .A3(new_n599), .A4(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n598), .A2(new_n527), .ZN(new_n1054));
  OAI21_X1  g629(.A(G1981), .B1(new_n1054), .B2(new_n595), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n993), .B2(new_n989), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1049), .A2(new_n1063), .A3(KEYINPUT52), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1049), .B2(KEYINPUT52), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1051), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1064), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1071), .A2(KEYINPUT114), .A3(new_n1051), .A4(new_n1062), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1038), .B(new_n1046), .C1(new_n1069), .C2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1006), .A2(new_n1009), .A3(new_n1024), .A4(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(G299), .B(KEYINPUT57), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NOR4_X1   g652(.A1(new_n959), .A2(new_n981), .A3(new_n965), .A4(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT115), .B(G1956), .Z(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1075), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1079), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n989), .A2(new_n1033), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n993), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n989), .A2(new_n991), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  XNOR2_X1  g662(.A(G299), .B(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n981), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n960), .A2(new_n1089), .A3(new_n993), .A4(new_n1076), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1081), .A2(KEYINPUT120), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n1075), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT121), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1092), .A2(new_n1098), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n987), .B2(new_n965), .ZN(new_n1105));
  NAND4_X1  g680(.A1(G160), .A2(new_n989), .A3(KEYINPUT116), .A4(G40), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT58), .B(G1341), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1103), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT118), .B(new_n1108), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n960), .A2(new_n1089), .A3(new_n993), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G1996), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1102), .B1(new_n1114), .B2(new_n623), .ZN(new_n1115));
  NAND2_X1  g690(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1107), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n564), .B(new_n1116), .C1(new_n1120), .C2(new_n1113), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1101), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT122), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1100), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1107), .A2(G2067), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n994), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n626), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n614), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1124), .A2(new_n1126), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1081), .B1(new_n1137), .B2(new_n626), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1091), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1074), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1020), .A2(new_n1141), .A3(new_n1023), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n1073), .A3(new_n1002), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1142), .A2(new_n1073), .A3(new_n1146), .A4(new_n1002), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1013), .A2(G8), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G286), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1073), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G1976), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1062), .A2(new_n1153), .A3(new_n771), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1053), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1060), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1046), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1067), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1045), .A2(G8), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1151), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1161), .A2(KEYINPUT63), .B1(new_n1158), .B2(new_n1046), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1152), .A2(new_n1156), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1148), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n978), .B1(new_n1140), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n967), .A2(new_n968), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n966), .B1(new_n1166), .B2(new_n818), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n966), .A2(new_n969), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1171));
  XNOR2_X1  g746(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n972), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n968), .B1(new_n1173), .B2(new_n971), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n966), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n966), .A2(new_n977), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  INV_X1    g752(.A(new_n966), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n974), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1172), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1165), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g756(.A(G229), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n878), .A2(new_n1183), .ZN(new_n1184));
  OR3_X1    g758(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1185));
  NOR3_X1   g759(.A1(new_n1184), .A2(new_n955), .A3(new_n1185), .ZN(G308));
  INV_X1    g760(.A(G308), .ZN(G225));
endmodule


