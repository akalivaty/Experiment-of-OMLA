

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  XOR2_X1 U325 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n294) );
  XNOR2_X1 U326 ( .A(G1GAT), .B(KEYINPUT104), .ZN(n293) );
  XNOR2_X1 U327 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U328 ( .A(KEYINPUT103), .B(n295), .Z(n457) );
  XOR2_X1 U329 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U330 ( .A(G141GAT), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U331 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U332 ( .A(G85GAT), .B(G162GAT), .Z(n299) );
  XNOR2_X1 U333 ( .A(G113GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U334 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U335 ( .A(n301), .B(n300), .ZN(n313) );
  XOR2_X1 U336 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n303) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n302) );
  XNOR2_X1 U338 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U339 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n305) );
  XNOR2_X1 U340 ( .A(KEYINPUT97), .B(G57GAT), .ZN(n304) );
  XNOR2_X1 U341 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U342 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U343 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n309) );
  XNOR2_X1 U344 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n308) );
  XNOR2_X1 U345 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U346 ( .A(KEYINPUT3), .B(n310), .ZN(n335) );
  XNOR2_X1 U347 ( .A(n311), .B(n335), .ZN(n312) );
  XNOR2_X1 U348 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(n314), .ZN(n320) );
  XOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT0), .Z(n316) );
  XNOR2_X1 U351 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n315) );
  XNOR2_X1 U352 ( .A(n316), .B(n315), .ZN(n345) );
  XOR2_X1 U353 ( .A(G134GAT), .B(n345), .Z(n318) );
  NAND2_X1 U354 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U355 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U356 ( .A(n320), .B(n319), .Z(n489) );
  INV_X1 U357 ( .A(n489), .ZN(n543) );
  XOR2_X1 U358 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n322) );
  XOR2_X1 U359 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n391) );
  XNOR2_X1 U361 ( .A(n431), .B(n391), .ZN(n321) );
  XNOR2_X1 U362 ( .A(n322), .B(n321), .ZN(n332) );
  XOR2_X1 U363 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n330) );
  XNOR2_X1 U364 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n323) );
  XNOR2_X1 U365 ( .A(n323), .B(KEYINPUT91), .ZN(n324) );
  XOR2_X1 U366 ( .A(n324), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U368 ( .A(n326), .B(n325), .ZN(n361) );
  XOR2_X1 U369 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U371 ( .A(n328), .B(n327), .ZN(n444) );
  XNOR2_X1 U372 ( .A(n361), .B(n444), .ZN(n329) );
  XNOR2_X1 U373 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U374 ( .A(n332), .B(n331), .Z(n334) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U376 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U377 ( .A(n336), .B(n335), .ZN(n545) );
  XOR2_X1 U378 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n338) );
  XNOR2_X1 U379 ( .A(KEYINPUT84), .B(KEYINPUT88), .ZN(n337) );
  XNOR2_X1 U380 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U381 ( .A(G176GAT), .B(KEYINPUT87), .Z(n340) );
  XOR2_X1 U382 ( .A(G113GAT), .B(G15GAT), .Z(n435) );
  XOR2_X1 U383 ( .A(G43GAT), .B(G134GAT), .Z(n395) );
  XNOR2_X1 U384 ( .A(n435), .B(n395), .ZN(n339) );
  XNOR2_X1 U385 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U386 ( .A(n342), .B(n341), .Z(n344) );
  NAND2_X1 U387 ( .A1(G227GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U388 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U389 ( .A(n346), .B(n345), .Z(n354) );
  XOR2_X1 U390 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n348) );
  XNOR2_X1 U391 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n347) );
  XNOR2_X1 U392 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U393 ( .A(n349), .B(KEYINPUT19), .Z(n351) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U395 ( .A(n351), .B(n350), .ZN(n365) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G71GAT), .ZN(n352) );
  XNOR2_X1 U397 ( .A(n352), .B(G120GAT), .ZN(n445) );
  XNOR2_X1 U398 ( .A(n365), .B(n445), .ZN(n353) );
  XOR2_X1 U399 ( .A(n354), .B(n353), .Z(n510) );
  INV_X1 U400 ( .A(n510), .ZN(n548) );
  XOR2_X1 U401 ( .A(G8GAT), .B(KEYINPUT77), .Z(n412) );
  XOR2_X1 U402 ( .A(n412), .B(KEYINPUT99), .Z(n356) );
  NAND2_X1 U403 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U404 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U405 ( .A(KEYINPUT100), .B(G92GAT), .Z(n358) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(G204GAT), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U408 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U409 ( .A(G176GAT), .B(G64GAT), .Z(n443) );
  XNOR2_X1 U410 ( .A(n361), .B(n443), .ZN(n362) );
  XNOR2_X1 U411 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U412 ( .A(n365), .B(n364), .ZN(n492) );
  INV_X1 U413 ( .A(n492), .ZN(n541) );
  NOR2_X1 U414 ( .A1(n548), .A2(n541), .ZN(n366) );
  NOR2_X1 U415 ( .A1(n545), .A2(n366), .ZN(n367) );
  XNOR2_X1 U416 ( .A(n367), .B(KEYINPUT25), .ZN(n370) );
  XNOR2_X1 U417 ( .A(n492), .B(KEYINPUT27), .ZN(n372) );
  NAND2_X1 U418 ( .A1(n545), .A2(n548), .ZN(n368) );
  XOR2_X1 U419 ( .A(n368), .B(KEYINPUT26), .Z(n564) );
  NAND2_X1 U420 ( .A1(n372), .A2(n564), .ZN(n369) );
  NAND2_X1 U421 ( .A1(n370), .A2(n369), .ZN(n371) );
  NAND2_X1 U422 ( .A1(n543), .A2(n371), .ZN(n376) );
  XOR2_X1 U423 ( .A(KEYINPUT89), .B(n548), .Z(n374) );
  XNOR2_X1 U424 ( .A(n545), .B(KEYINPUT28), .ZN(n513) );
  NAND2_X1 U425 ( .A1(n489), .A2(n372), .ZN(n509) );
  NOR2_X1 U426 ( .A1(n513), .A2(n509), .ZN(n373) );
  NAND2_X1 U427 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U428 ( .A1(n376), .A2(n375), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n377), .B(KEYINPUT101), .ZN(n464) );
  XOR2_X1 U430 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n379) );
  XNOR2_X1 U431 ( .A(G36GAT), .B(G29GAT), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(n380), .Z(n440) );
  INV_X1 U434 ( .A(n440), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT11), .B(G106GAT), .Z(n382) );
  XNOR2_X1 U436 ( .A(G190GAT), .B(G99GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n399) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n386) );
  XNOR2_X1 U440 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT75), .Z(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U445 ( .A(n390), .B(n389), .Z(n397) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G92GAT), .Z(n451) );
  XOR2_X1 U447 ( .A(n451), .B(n391), .Z(n393) );
  NAND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U452 ( .A(n399), .B(n398), .Z(n559) );
  XOR2_X1 U453 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n401) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G64GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n419) );
  XOR2_X1 U460 ( .A(G127GAT), .B(G71GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(G15GAT), .B(G183GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U463 ( .A(G78GAT), .B(G211GAT), .Z(n409) );
  XNOR2_X1 U464 ( .A(G22GAT), .B(G155GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U466 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U467 ( .A(G57GAT), .B(KEYINPUT13), .Z(n442) );
  XOR2_X1 U468 ( .A(KEYINPUT81), .B(n412), .Z(n414) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n442), .B(n415), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U473 ( .A(n419), .B(n418), .Z(n577) );
  NOR2_X1 U474 ( .A1(n559), .A2(n577), .ZN(n420) );
  XOR2_X1 U475 ( .A(KEYINPUT16), .B(n420), .Z(n421) );
  NOR2_X1 U476 ( .A1(n464), .A2(n421), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT102), .B(n422), .Z(n478) );
  XOR2_X1 U478 ( .A(KEYINPUT70), .B(KEYINPUT66), .Z(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n439) );
  XOR2_X1 U481 ( .A(G197GAT), .B(G50GAT), .Z(n426) );
  XNOR2_X1 U482 ( .A(G169GAT), .B(G43GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U484 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n428) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n437) );
  XOR2_X1 U488 ( .A(n431), .B(G8GAT), .Z(n433) );
  NAND2_X1 U489 ( .A1(G229GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n550) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n455) );
  XOR2_X1 U498 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n449) );
  XNOR2_X1 U499 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U501 ( .A(n451), .B(n450), .Z(n453) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n573) );
  NAND2_X1 U505 ( .A1(n550), .A2(n573), .ZN(n467) );
  NOR2_X1 U506 ( .A1(n478), .A2(n467), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n462), .A2(n489), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n457), .B(n456), .ZN(G1324GAT) );
  NAND2_X1 U509 ( .A1(n492), .A2(n462), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n458), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n460) );
  NAND2_X1 U512 ( .A1(n462), .A2(n510), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(G15GAT), .B(n461), .ZN(G1326GAT) );
  NAND2_X1 U515 ( .A1(n513), .A2(n462), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U517 ( .A(G29GAT), .B(KEYINPUT39), .Z(n471) );
  XOR2_X1 U518 ( .A(KEYINPUT36), .B(n559), .Z(n581) );
  NOR2_X1 U519 ( .A1(n464), .A2(n581), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n577), .ZN(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT37), .B(n466), .Z(n486) );
  NOR2_X1 U522 ( .A1(n486), .A2(n467), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n468) );
  XNOR2_X1 U524 ( .A(n469), .B(n468), .ZN(n475) );
  NAND2_X1 U525 ( .A1(n489), .A2(n475), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(G1328GAT) );
  NAND2_X1 U527 ( .A1(n475), .A2(n492), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U529 ( .A1(n475), .A2(n510), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT40), .ZN(n474) );
  XNOR2_X1 U531 ( .A(G43GAT), .B(n474), .ZN(G1330GAT) );
  NAND2_X1 U532 ( .A1(n475), .A2(n513), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U534 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n480) );
  XOR2_X1 U535 ( .A(n573), .B(KEYINPUT41), .Z(n529) );
  INV_X1 U536 ( .A(n529), .ZN(n553) );
  INV_X1 U537 ( .A(n550), .ZN(n568) );
  NAND2_X1 U538 ( .A1(n553), .A2(n568), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(KEYINPUT108), .ZN(n487) );
  NOR2_X1 U540 ( .A1(n487), .A2(n478), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n489), .A2(n483), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(G1332GAT) );
  NAND2_X1 U543 ( .A1(n492), .A2(n483), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U545 ( .A1(n510), .A2(n483), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n482), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U547 ( .A(G78GAT), .B(KEYINPUT43), .Z(n485) );
  NAND2_X1 U548 ( .A1(n483), .A2(n513), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(G1335GAT) );
  NOR2_X1 U550 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U551 ( .A(KEYINPUT109), .B(n488), .Z(n495) );
  NAND2_X1 U552 ( .A1(n495), .A2(n489), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT110), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(n491), .ZN(G1336GAT) );
  NAND2_X1 U555 ( .A1(n492), .A2(n495), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U557 ( .A1(n510), .A2(n495), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U559 ( .A1(n513), .A2(n495), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT44), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G106GAT), .B(n497), .ZN(G1339GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n515) );
  INV_X1 U563 ( .A(n559), .ZN(n538) );
  INV_X1 U564 ( .A(n577), .ZN(n557) );
  NOR2_X1 U565 ( .A1(n568), .A2(n529), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n498), .B(KEYINPUT46), .ZN(n499) );
  NOR2_X1 U567 ( .A1(n557), .A2(n499), .ZN(n500) );
  NAND2_X1 U568 ( .A1(n538), .A2(n500), .ZN(n501) );
  XNOR2_X1 U569 ( .A(KEYINPUT47), .B(n501), .ZN(n507) );
  NOR2_X1 U570 ( .A1(n581), .A2(n577), .ZN(n503) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n503), .B(n502), .ZN(n505) );
  NAND2_X1 U573 ( .A1(n568), .A2(n573), .ZN(n504) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n506) );
  NOR2_X1 U575 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT48), .ZN(n540) );
  NOR2_X1 U577 ( .A1(n540), .A2(n509), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n526), .A2(n510), .ZN(n511) );
  XOR2_X1 U579 ( .A(KEYINPUT111), .B(n511), .Z(n512) );
  NOR2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n550), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G113GAT), .B(n516), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U585 ( .A1(n522), .A2(n553), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n520) );
  NAND2_X1 U588 ( .A1(n522), .A2(n557), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U590 ( .A(G127GAT), .B(n521), .Z(G1342GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U592 ( .A1(n522), .A2(n559), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U594 ( .A(G134GAT), .B(n525), .Z(G1343GAT) );
  NAND2_X1 U595 ( .A1(n526), .A2(n564), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n568), .A2(n537), .ZN(n527) );
  XOR2_X1 U597 ( .A(G141GAT), .B(n527), .Z(n528) );
  XNOR2_X1 U598 ( .A(KEYINPUT116), .B(n528), .ZN(G1344GAT) );
  NOR2_X1 U599 ( .A1(n529), .A2(n537), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n531) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n530) );
  XNOR2_X1 U602 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U603 ( .A(KEYINPUT52), .B(n532), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n577), .A2(n537), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(G1346GAT) );
  NOR2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U609 ( .A(G162GAT), .B(n539), .Z(G1347GAT) );
  XOR2_X1 U610 ( .A(G169GAT), .B(KEYINPUT121), .Z(n552) );
  NOR2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n542), .B(KEYINPUT54), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n565) );
  NOR2_X1 U614 ( .A1(n545), .A2(n565), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n546), .B(KEYINPUT55), .ZN(n547) );
  NOR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(KEYINPUT120), .B(n549), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n560), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G190GAT), .B(n563), .Z(G1351GAT) );
  INV_X1 U630 ( .A(n564), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT123), .B(n567), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n568), .A2(n580), .ZN(n572) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT124), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n580), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n578), .Z(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

