//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AND2_X1   g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G87), .C2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G50), .A2(G226), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n233), .A2(G50), .A3(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n213), .B(new_n229), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n218), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT67), .B(G250), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n230), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n254), .B2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT8), .B(G58), .Z(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(new_n264), .B1(G150), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT68), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n259), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n269), .B2(new_n259), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n257), .B(new_n261), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G222), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G223), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(G77), .C2(new_n275), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(G1), .B(G13), .C1(new_n263), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n281), .B(new_n284), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n289), .A2(G179), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n274), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(new_n254), .A3(G13), .A4(G20), .ZN(new_n296));
  AOI21_X1  g0096(.A(G77), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n260), .A2(new_n295), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n215), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n262), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n300));
  INV_X1    g0100(.A(new_n264), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT15), .B(G87), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g0103(.A(new_n297), .B(new_n299), .C1(new_n259), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n284), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n275), .A2(G232), .A3(new_n277), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n307));
  INV_X1    g0107(.A(G107), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n275), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n305), .B1(new_n309), .B2(new_n280), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n287), .A2(G244), .A3(new_n282), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT72), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n304), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n290), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n274), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n273), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n271), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n324), .A2(KEYINPUT9), .A3(new_n257), .A4(new_n261), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT71), .B(G200), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n289), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n289), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n322), .A2(new_n325), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n293), .B(new_n320), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  INV_X1    g0135(.A(new_n262), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n255), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n260), .B2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n275), .B2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT76), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n231), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n339), .ZN(new_n349));
  OAI21_X1  g0149(.A(G68), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n225), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n265), .A2(G159), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT16), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n344), .B2(new_n231), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n339), .B(G20), .C1(new_n341), .C2(new_n343), .ZN(new_n359));
  OAI21_X1  g0159(.A(G68), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n259), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n338), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT77), .B(new_n338), .C1(new_n357), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G232), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n284), .B1(new_n288), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n285), .A2(G1698), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n275), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n280), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n284), .B(KEYINPUT78), .C1(new_n288), .C2(new_n368), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n371), .A2(new_n377), .A3(new_n311), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n287), .B1(new_n374), .B2(new_n375), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n290), .B1(new_n380), .B2(new_n369), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n335), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g0184(.A(KEYINPUT18), .B(new_n382), .C1(new_n365), .C2(new_n366), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n341), .A2(new_n343), .A3(G232), .A4(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n275), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n275), .A2(G226), .A3(new_n277), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n280), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n284), .B1(new_n288), .B2(new_n226), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n387), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI211_X1 g0198(.A(KEYINPUT13), .B(new_n396), .C1(new_n394), .C2(new_n280), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n397), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT13), .ZN(new_n403));
  OAI21_X1  g0203(.A(G179), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n398), .B2(new_n399), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(G169), .C1(new_n398), .C2(new_n399), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT12), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n410), .B(G68), .C1(new_n294), .C2(new_n296), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n225), .B1(new_n298), .B2(KEYINPUT12), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n410), .C2(new_n255), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n265), .A2(G50), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT75), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n415), .B1(new_n231), .B2(G68), .C1(new_n215), .C2(new_n301), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n416), .A2(new_n417), .A3(new_n259), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n416), .B2(new_n259), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n401), .A2(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n395), .A2(new_n387), .A3(new_n397), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n402), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n399), .B1(new_n398), .B2(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n420), .B1(new_n425), .B2(G190), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n398), .B2(new_n399), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n409), .A2(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n371), .A2(new_n377), .A3(new_n329), .A4(new_n378), .ZN(new_n429));
  INV_X1    g0229(.A(G200), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n380), .B2(new_n369), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n338), .B(new_n432), .C1(new_n357), .C2(new_n362), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT17), .B1(new_n433), .B2(KEYINPUT79), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT79), .B1(new_n433), .B2(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT79), .B(KEYINPUT17), .C1(new_n433), .C2(KEYINPUT80), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n318), .A2(new_n327), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n304), .B(new_n439), .C1(new_n329), .C2(new_n318), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n386), .A2(new_n428), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n334), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n254), .A2(G33), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(new_n258), .A3(G116), .A4(new_n230), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n444), .A2(new_n294), .A3(new_n296), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n294), .B2(new_n296), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n258), .A2(new_n230), .B1(G20), .B2(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n231), .C1(G33), .C2(new_n217), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n448), .A2(KEYINPUT20), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT20), .B1(new_n448), .B2(new_n450), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n445), .A2(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n254), .A2(G45), .A3(G274), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n254), .A2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n280), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n462), .B2(G270), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n341), .A2(new_n343), .A3(G257), .A4(new_n277), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n341), .A2(new_n343), .A3(G264), .A4(G1698), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n275), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n280), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n468), .A3(G190), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n463), .A2(new_n468), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n454), .B(new_n469), .C1(new_n470), .C2(new_n430), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n463), .A2(new_n468), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G169), .A3(new_n453), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT21), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(G179), .A3(new_n453), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n290), .B1(new_n463), .B2(new_n468), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT21), .A3(new_n453), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n471), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT84), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n341), .A2(new_n343), .A3(G244), .A4(new_n277), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n275), .A2(G244), .A3(new_n485), .A4(new_n277), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n486), .A3(new_n449), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n280), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n459), .B1(new_n462), .B2(G257), .ZN(new_n490));
  AOI21_X1  g0290(.A(G169), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(G107), .B1(new_n346), .B2(new_n349), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n265), .A2(G77), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n308), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  XOR2_X1   g0294(.A(G97), .B(G107), .Z(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n259), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n255), .A2(G97), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n255), .A2(new_n443), .A3(new_n230), .A4(new_n258), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n217), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n491), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n489), .A2(new_n490), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G179), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n259), .ZN(new_n509));
  NAND3_X1  g0309(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n231), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n217), .A3(new_n308), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n231), .A2(G33), .A3(G97), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n511), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n341), .A2(new_n343), .A3(new_n231), .A4(G68), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT15), .B(G87), .Z(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n294), .B2(new_n296), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n501), .A2(new_n512), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n226), .A2(new_n277), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n216), .A2(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n341), .A2(new_n523), .A3(new_n343), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n280), .ZN(new_n528));
  XOR2_X1   g0328(.A(new_n456), .B(KEYINPUT83), .Z(new_n529));
  NAND3_X1  g0329(.A1(new_n287), .A2(G250), .A3(new_n460), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(G190), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n287), .B1(new_n525), .B2(new_n526), .ZN(new_n532));
  INV_X1    g0332(.A(new_n530), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n456), .B(KEYINPUT83), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n522), .B(new_n531), .C1(new_n535), .C2(new_n326), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n511), .A2(new_n513), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n514), .A2(new_n515), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n517), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n259), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n501), .A2(new_n302), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n294), .A2(new_n296), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n302), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n528), .A2(new_n311), .A3(new_n529), .A4(new_n530), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n535), .C2(G169), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n341), .A2(new_n343), .A3(new_n231), .A4(G87), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n275), .A2(KEYINPUT22), .A3(new_n231), .A4(G87), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n231), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n308), .A2(KEYINPUT23), .A3(G20), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n554), .B1(new_n264), .B2(G116), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT24), .A4(new_n555), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n259), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n501), .A2(new_n308), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n255), .A2(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT25), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n341), .A2(new_n343), .A3(G257), .A4(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n341), .A2(new_n343), .A3(G250), .A4(new_n277), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n566), .C1(new_n263), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n280), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n462), .A2(G264), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n311), .A2(new_n569), .A3(new_n458), .A4(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n568), .A2(new_n280), .B1(new_n462), .B2(G264), .ZN(new_n572));
  AOI21_X1  g0372(.A(G169), .B1(new_n572), .B2(new_n458), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n547), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n502), .B1(new_n498), .B2(new_n259), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT82), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n489), .A2(new_n577), .A3(G190), .A4(new_n490), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n505), .A2(G200), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT82), .B1(new_n505), .B2(new_n329), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n569), .A2(new_n570), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n459), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G190), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n582), .B(new_n585), .C1(new_n430), .C2(new_n584), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n508), .A2(new_n575), .A3(new_n581), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n481), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n442), .A2(new_n588), .ZN(G372));
  INV_X1    g0389(.A(new_n293), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n332), .A2(new_n333), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n363), .A2(new_n383), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(new_n335), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n426), .A2(new_n427), .ZN(new_n595));
  INV_X1    g0395(.A(new_n320), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n406), .A2(new_n408), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n311), .B1(new_n423), .B2(new_n424), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n420), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n601), .B2(new_n438), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(KEYINPUT86), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n602), .A2(KEYINPUT86), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n590), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n477), .A2(KEYINPUT21), .A3(new_n453), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT21), .B1(new_n477), .B2(new_n453), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n574), .A2(new_n564), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n476), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n547), .A2(KEYINPUT85), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n536), .A2(new_n546), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n614), .A3(new_n586), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n508), .A2(new_n581), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n546), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n576), .A2(new_n491), .A3(new_n506), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT26), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n547), .ZN(new_n620));
  AND4_X1   g0420(.A1(KEYINPUT26), .A2(new_n504), .A3(new_n620), .A4(new_n507), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n442), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n605), .A2(new_n623), .ZN(G369));
  NOR2_X1   g0424(.A1(new_n209), .A2(G20), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OR3_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .A3(G1), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT27), .B1(new_n626), .B2(G1), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n609), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n564), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n586), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n609), .ZN(new_n635));
  INV_X1    g0435(.A(new_n632), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n608), .A2(new_n476), .ZN(new_n641));
  INV_X1    g0441(.A(new_n631), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n632), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n642), .A2(new_n454), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n481), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n640), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n651), .ZN(G399));
  INV_X1    g0452(.A(new_n211), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G41), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n254), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n513), .A2(G116), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n655), .A2(new_n656), .B1(new_n236), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT28), .Z(new_n658));
  NOR2_X1   g0458(.A1(new_n617), .A2(new_n622), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n631), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT29), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n504), .A2(new_n620), .A3(new_n507), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n662), .A2(KEYINPUT89), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT89), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n614), .A2(KEYINPUT26), .A3(new_n618), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(KEYINPUT29), .B(new_n642), .C1(new_n667), .C2(new_n617), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n584), .A2(new_n470), .ZN(new_n670));
  INV_X1    g0470(.A(new_n535), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n311), .A3(new_n671), .A4(new_n505), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n463), .A2(new_n468), .A3(G179), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n505), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n535), .A2(new_n572), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NOR4_X1   g0478(.A1(new_n505), .A2(new_n676), .A3(new_n674), .A4(KEYINPUT30), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n672), .B(KEYINPUT88), .C1(new_n678), .C2(new_n679), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n631), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n588), .A2(new_n642), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n669), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n658), .B1(new_n691), .B2(G1), .ZN(G364));
  AOI21_X1  g0492(.A(new_n254), .B1(new_n625), .B2(G45), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n654), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n650), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(G330), .B2(new_n648), .ZN(new_n697));
  INV_X1    g0497(.A(new_n695), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n326), .A2(G179), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n231), .A2(G190), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(G20), .A3(G190), .ZN(new_n703));
  OAI221_X1 g0503(.A(new_n275), .B1(new_n702), .B2(new_n308), .C1(new_n512), .C2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n430), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(G50), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(G20), .A2(G179), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n708), .A2(G190), .A3(G200), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n215), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G179), .A2(G200), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G159), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT32), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n705), .A2(G200), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n231), .B1(new_n712), .B2(G190), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n708), .A2(new_n430), .A3(G190), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n720), .A2(G97), .B1(G68), .B2(new_n721), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n716), .B1(new_n718), .B2(new_n351), .C1(new_n722), .C2(KEYINPUT92), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n711), .B(new_n723), .C1(KEYINPUT92), .C2(new_n722), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n707), .B(new_n724), .C1(KEYINPUT32), .C2(new_n715), .ZN(new_n725));
  INV_X1    g0525(.A(new_n706), .ZN(new_n726));
  INV_X1    g0526(.A(G326), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G311), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n710), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G329), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n344), .B1(new_n719), .B2(new_n567), .C1(new_n731), .C2(new_n713), .ZN(new_n732));
  INV_X1    g0532(.A(new_n702), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n730), .B(new_n732), .C1(new_n733), .C2(G283), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(G317), .ZN(new_n736));
  INV_X1    g0536(.A(new_n721), .ZN(new_n737));
  INV_X1    g0537(.A(G322), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n736), .A2(new_n737), .B1(new_n718), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n734), .B(new_n740), .C1(new_n466), .C2(new_n703), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n725), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n230), .B1(G20), .B2(new_n290), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(G355), .A2(new_n211), .A3(new_n275), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n249), .A2(G45), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT90), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n653), .A2(new_n275), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n235), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n745), .B1(G116), .B2(new_n211), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n647), .B(new_n751), .C1(new_n481), .C2(new_n646), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n744), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n697), .B1(new_n698), .B2(new_n755), .ZN(G396));
  AND3_X1   g0556(.A1(new_n317), .A2(new_n319), .A3(new_n642), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n304), .A2(new_n642), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n317), .A2(new_n319), .B1(new_n440), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n660), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n689), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT96), .Z(new_n763));
  AOI21_X1  g0563(.A(new_n695), .B1(new_n761), .B2(new_n689), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n760), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n733), .A2(G87), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n720), .A2(G97), .B1(G294), .B2(new_n717), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n344), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n703), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G116), .A2(new_n709), .B1(new_n706), .B2(G303), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(new_n737), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT95), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n772), .A2(G107), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n771), .B(new_n778), .C1(G311), .C2(new_n714), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n733), .A2(G68), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G159), .A2(new_n709), .B1(new_n717), .B2(G143), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n706), .A2(G137), .ZN(new_n782));
  INV_X1    g0582(.A(G150), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n737), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT34), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(new_n785), .B1(G132), .B2(new_n714), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n720), .A2(G58), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n780), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n344), .B(new_n789), .C1(G50), .C2(new_n772), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n743), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n743), .A2(new_n767), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n215), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n768), .A2(new_n695), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n765), .A2(new_n794), .ZN(G384));
  NAND2_X1  g0595(.A1(new_n684), .A2(new_n685), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n479), .B(KEYINPUT84), .ZN(new_n797));
  INV_X1    g0597(.A(new_n616), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n575), .A2(new_n586), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n642), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n631), .A4(new_n683), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n760), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n420), .A2(new_n631), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n595), .A2(new_n600), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT98), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n595), .A2(new_n600), .A3(KEYINPUT98), .A4(new_n804), .ZN(new_n808));
  INV_X1    g0608(.A(new_n600), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n807), .A2(new_n808), .B1(new_n809), .B2(new_n631), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT38), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n225), .B1(new_n340), .B2(new_n345), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n355), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n509), .B1(new_n814), .B2(KEYINPUT16), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n347), .B1(new_n358), .B2(new_n359), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n355), .B1(new_n818), .B2(G68), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n815), .B1(new_n819), .B2(KEYINPUT16), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT77), .B1(new_n820), .B2(new_n338), .ZN(new_n821));
  INV_X1    g0621(.A(new_n366), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n383), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n629), .B(KEYINPUT100), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n821), .B2(new_n822), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n826), .A3(new_n827), .A4(new_n433), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT16), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n813), .B2(new_n355), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n361), .A2(new_n830), .A3(new_n259), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n338), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n383), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT99), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n433), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n629), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n834), .B1(new_n833), .B2(new_n433), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n823), .A2(KEYINPUT18), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n367), .A2(new_n335), .A3(new_n383), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n438), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n837), .ZN(new_n844));
  AOI221_X4 g0644(.A(new_n812), .B1(new_n828), .B2(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n438), .A2(new_n593), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n824), .B1(new_n365), .B2(new_n366), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n433), .ZN(new_n849));
  INV_X1    g0649(.A(new_n592), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n828), .B1(new_n851), .B2(new_n827), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n811), .B(KEYINPUT40), .C1(new_n845), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n837), .B1(new_n386), .B2(new_n438), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n828), .A2(new_n840), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n812), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n843), .A2(new_n844), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n828), .A2(new_n840), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n855), .B(KEYINPUT40), .C1(new_n811), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n766), .B1(new_n686), .B2(new_n801), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n809), .A2(new_n631), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT98), .B1(new_n428), .B2(new_n804), .ZN(new_n866));
  INV_X1    g0666(.A(new_n808), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n859), .B2(new_n860), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n864), .B(new_n868), .C1(new_n845), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT101), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(G330), .B(new_n854), .C1(new_n863), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n442), .A2(G330), .A3(new_n802), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n845), .A2(new_n869), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n868), .A2(new_n760), .A3(new_n802), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n855), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n870), .A2(KEYINPUT101), .A3(new_n871), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n881), .A2(new_n442), .A3(new_n802), .A4(new_n854), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n593), .A2(new_n825), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n642), .B(new_n760), .C1(new_n617), .C2(new_n622), .ZN(new_n885));
  INV_X1    g0685(.A(new_n757), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n876), .A2(new_n810), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n809), .A2(new_n642), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n845), .B2(new_n853), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n858), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n884), .B(new_n889), .C1(new_n891), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n883), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n442), .A2(new_n668), .A3(new_n661), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n605), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n254), .B2(new_n625), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n496), .B(KEYINPUT97), .Z(new_n903));
  AOI21_X1  g0703(.A(new_n446), .B1(new_n903), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n232), .C1(KEYINPUT35), .C2(new_n903), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n235), .A2(new_n215), .A3(new_n352), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n225), .A2(G50), .ZN(new_n908));
  OAI211_X1 g0708(.A(G1), .B(new_n209), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(new_n906), .A3(new_n909), .ZN(G367));
  INV_X1    g0710(.A(new_n640), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n643), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n637), .A2(KEYINPUT87), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n644), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n649), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n650), .A3(new_n915), .ZN(new_n918));
  AND4_X1   g0718(.A1(new_n689), .A2(new_n917), .A3(new_n669), .A4(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n636), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n798), .B1(new_n576), .B2(new_n642), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n618), .A2(new_n631), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n645), .A2(new_n925), .A3(new_n920), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT44), .B1(new_n645), .B2(new_n925), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT44), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n929), .A2(new_n651), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n930), .A2(new_n927), .A3(new_n928), .A4(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n650), .A3(new_n640), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n919), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT107), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n919), .A2(new_n933), .A3(new_n935), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n690), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n654), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n693), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT42), .B1(new_n915), .B2(new_n926), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n508), .B1(new_n923), .B2(new_n609), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n642), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT42), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n640), .A2(new_n947), .A3(new_n644), .A4(new_n925), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n642), .A2(new_n522), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n614), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n951), .A2(new_n546), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT102), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n949), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT105), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n958), .B2(new_n949), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT103), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT104), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n651), .A2(new_n926), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n961), .B(KEYINPUT103), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(KEYINPUT104), .A3(new_n960), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n968), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n969), .A2(KEYINPUT104), .A3(new_n960), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT104), .B1(new_n969), .B2(new_n960), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n943), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n733), .A2(G77), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n719), .A2(new_n225), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G150), .B2(new_n717), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n344), .B(new_n982), .C1(G143), .C2(new_n706), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n772), .A2(G58), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G50), .A2(new_n709), .B1(new_n721), .B2(G159), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT109), .B(G137), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n714), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n702), .A2(new_n217), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G303), .B2(new_n717), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n774), .B2(new_n710), .C1(new_n729), .C2(new_n726), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G317), .B2(new_n714), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n772), .A2(G116), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n275), .B1(new_n720), .B2(G107), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n737), .A2(new_n567), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n988), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n743), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n954), .A2(new_n751), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n748), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n752), .B1(new_n211), .B2(new_n302), .C1(new_n245), .C2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n695), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n976), .A2(new_n1004), .ZN(G387));
  AOI21_X1  g0805(.A(new_n698), .B1(new_n911), .B2(new_n751), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n653), .A2(G107), .ZN(new_n1007));
  INV_X1    g0807(.A(G45), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n241), .A2(new_n1008), .A3(new_n275), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n336), .A2(G50), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT50), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1010), .A2(new_n1013), .B1(new_n225), .B2(new_n215), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n344), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n656), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n752), .B(new_n1007), .C1(new_n1016), .C2(new_n653), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(G159), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n726), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n719), .A2(new_n302), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n989), .B1(G150), .B2(new_n714), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n772), .A2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n275), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT110), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1020), .B(new_n1021), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n717), .A2(G50), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n262), .A2(new_n721), .B1(new_n709), .B2(G68), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G311), .A2(new_n721), .B1(new_n706), .B2(G322), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n466), .B2(new_n710), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G317), .B2(new_n717), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT48), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n774), .B2(new_n719), .C1(new_n567), .C2(new_n703), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT49), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n344), .B1(new_n727), .B2(new_n713), .C1(new_n702), .C2(new_n446), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n743), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n917), .A2(new_n918), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n694), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n654), .B1(new_n1041), .B2(new_n691), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n919), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n937), .A2(new_n939), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n933), .A2(new_n935), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n654), .C1(new_n1046), .C2(new_n919), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n694), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n926), .A2(new_n751), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT112), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n752), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n211), .A2(new_n217), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n748), .C2(new_n252), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n772), .A2(G68), .B1(G143), .B2(new_n714), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT113), .ZN(new_n1055));
  INV_X1    g0855(.A(G50), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n275), .B1(new_n737), .B2(new_n1056), .C1(new_n336), .C2(new_n710), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G77), .B2(new_n720), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G150), .A2(new_n706), .B1(new_n717), .B2(G159), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT51), .Z(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n769), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n703), .A2(new_n774), .B1(new_n702), .B2(new_n308), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n717), .B1(new_n706), .B2(G317), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n275), .B1(G294), .B2(new_n709), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n446), .B2(new_n719), .C1(new_n738), .C2(new_n713), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n466), .B2(new_n737), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1061), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n698), .B(new_n1053), .C1(new_n1069), .C2(new_n743), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1050), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1047), .A2(new_n1048), .A3(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n895), .A2(new_n767), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n344), .B1(new_n733), .B2(G50), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT54), .B(G143), .Z(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n709), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n721), .A2(new_n986), .B1(new_n706), .B2(G128), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G125), .A2(new_n714), .B1(new_n720), .B2(G159), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n703), .A2(new_n783), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1081), .B(new_n1085), .C1(G132), .C2(new_n717), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n780), .B1(new_n512), .B2(new_n703), .C1(new_n774), .C2(new_n726), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n710), .A2(new_n217), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n344), .B1(new_n719), .B2(new_n215), .C1(new_n567), .C2(new_n713), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n737), .A2(new_n308), .B1(new_n718), .B2(new_n446), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n743), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n792), .A2(new_n336), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1073), .A2(new_n695), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n811), .A2(G330), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n891), .B1(new_n868), .B2(new_n887), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n893), .B2(new_n894), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n890), .B1(new_n845), .B2(new_n853), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n759), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n642), .B(new_n1101), .C1(new_n667), .C2(new_n617), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n810), .B1(new_n886), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1095), .B(new_n1097), .C1(new_n1099), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n868), .A2(new_n688), .A3(G330), .A4(new_n760), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1095), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1097), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT115), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n693), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1108), .B(new_n1114), .C1(new_n896), .C2(new_n1098), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1105), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT115), .B1(new_n1117), .B2(new_n694), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1094), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n605), .A2(new_n899), .A3(new_n874), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1102), .A2(new_n886), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(G330), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n810), .B1(new_n803), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1108), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n810), .B1(new_n689), .B2(new_n766), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n888), .B1(new_n1126), .B2(new_n1096), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1116), .B2(new_n1105), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1111), .A2(new_n1128), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n654), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1119), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(G378));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n331), .B(KEYINPUT10), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n274), .A2(new_n836), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n293), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1137), .B2(new_n293), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1139), .A3(new_n1135), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n873), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n881), .A2(G330), .A3(new_n854), .A4(new_n1145), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1147), .A2(new_n1148), .A3(new_n897), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n897), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n605), .A2(new_n899), .A3(new_n874), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1149), .A2(new_n1150), .B1(new_n1129), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n654), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1152), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1111), .B2(new_n1128), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(KEYINPUT57), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n654), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n694), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1146), .A2(new_n767), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n772), .A2(new_n1077), .B1(G137), .B2(new_n709), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G132), .A2(new_n721), .B1(new_n706), .B2(G125), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n783), .C2(new_n719), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G128), .B2(new_n717), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT59), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n714), .C2(G124), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n1019), .C2(new_n702), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n978), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n286), .B(new_n344), .C1(new_n737), .C2(new_n217), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n733), .B2(G58), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n446), .B2(new_n726), .C1(new_n774), .C2(new_n713), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n519), .B2(new_n709), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n717), .A2(G107), .ZN(new_n1178));
  AND4_X1   g0978(.A1(new_n1173), .A2(new_n1177), .A3(new_n1023), .A4(new_n1178), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G50), .B1(new_n344), .B2(new_n286), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(G33), .B2(G41), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT118), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1172), .A2(new_n1180), .A3(new_n1181), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n743), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n792), .A2(new_n1056), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1165), .A2(new_n695), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1164), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1163), .A2(new_n1192), .ZN(G375));
  NOR2_X1   g0993(.A1(new_n1127), .A2(new_n1125), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n693), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n733), .A2(G58), .B1(G128), .B2(new_n714), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n706), .A2(G132), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1196), .B1(KEYINPUT121), .B2(new_n1197), .C1(new_n783), .C2(new_n710), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(KEYINPUT121), .B2(new_n1197), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n772), .A2(G159), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n720), .A2(G50), .B1(new_n1077), .B2(new_n721), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n344), .B1(new_n717), .B2(new_n986), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n977), .B1(new_n217), .B2(new_n703), .C1(new_n774), .C2(new_n718), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1021), .B(new_n1204), .C1(G107), .C2(new_n709), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G116), .A2(new_n721), .B1(new_n706), .B2(G294), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n344), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n713), .A2(new_n466), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1203), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT122), .Z(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n743), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n792), .A2(new_n225), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n810), .A2(new_n767), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n695), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1195), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1194), .A2(new_n1151), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1128), .A2(new_n1217), .A3(new_n941), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(G381));
  NOR2_X1   g1019(.A1(G375), .A2(G378), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1004), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n973), .A2(new_n974), .A3(new_n972), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n968), .B1(new_n967), .B2(new_n970), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1221), .B1(new_n1224), .B2(new_n943), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  OR3_X1    g1026(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G396), .A2(new_n1226), .A3(G393), .A4(new_n1227), .ZN(G407));
  INV_X1    g1028(.A(G213), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(G343), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT124), .Z(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1220), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G407), .A2(new_n1232), .ZN(G409));
  NAND3_X1  g1033(.A1(new_n976), .A2(new_n1004), .A3(G390), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(G393), .B(G396), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1235), .B(G390), .C1(new_n976), .C2(new_n1004), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(KEYINPUT126), .ZN(new_n1237));
  INV_X1    g1037(.A(G390), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(G387), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1234), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1237), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1234), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n654), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n654), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1158), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(G378), .B1(new_n1250), .B2(new_n1191), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1230), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1192), .B1(new_n942), .B2(new_n1153), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G378), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1217), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1194), .A2(KEYINPUT60), .A3(new_n1151), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n654), .A3(new_n1128), .A4(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1216), .A2(G384), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1216), .B2(new_n1259), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1251), .A2(new_n1252), .A3(new_n1255), .A4(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1133), .B1(new_n1163), .B2(new_n1192), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1265), .A2(new_n1231), .A3(new_n1254), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1263), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n1246), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1246), .A2(new_n1264), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1230), .A2(G2897), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G2897), .B(new_n1231), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G2897), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1216), .A2(new_n1259), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1279), .B2(new_n1260), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1231), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1272), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1270), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1245), .B1(new_n1269), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1267), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1251), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1280), .A2(KEYINPUT125), .A3(new_n1231), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1289), .A2(new_n1290), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1285), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1264), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1244), .B(new_n1287), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(new_n1294), .ZN(G405));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1234), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1241), .B1(new_n1225), .B2(G390), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1235), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G387), .A2(new_n1238), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1301), .B2(new_n1242), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1240), .A2(KEYINPUT127), .A3(new_n1243), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  OR3_X1    g1104(.A1(new_n1220), .A2(new_n1265), .A3(new_n1263), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1263), .B1(new_n1220), .B2(new_n1265), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1305), .A2(new_n1306), .B1(new_n1296), .B2(new_n1244), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(G402));
endmodule


