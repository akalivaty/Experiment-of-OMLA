

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n701), .B(KEYINPUT64), .ZN(n706) );
  BUF_X1 U553 ( .A(n579), .Z(n561) );
  BUF_X1 U554 ( .A(n571), .Z(n562) );
  NAND2_X2 U555 ( .A1(n754), .A2(G8), .ZN(n789) );
  XNOR2_X1 U556 ( .A(n523), .B(n522), .ZN(n571) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NAND2_X1 U558 ( .A1(n571), .A2(G137), .ZN(n572) );
  XNOR2_X1 U559 ( .A(n706), .B(n705), .ZN(n736) );
  NOR2_X1 U560 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U561 ( .A(n735), .B(n734), .ZN(n742) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n789), .ZN(n766) );
  INV_X1 U563 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U564 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U565 ( .A1(n574), .A2(KEYINPUT69), .ZN(n575) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n526), .ZN(n559) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(n774), .Z(n519) );
  NOR2_X2 U568 ( .A1(n583), .A2(n582), .ZN(G160) );
  INV_X1 U569 ( .A(KEYINPUT94), .ZN(n705) );
  INV_X1 U570 ( .A(KEYINPUT28), .ZN(n710) );
  INV_X1 U571 ( .A(KEYINPUT29), .ZN(n734) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n522) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  AND2_X1 U574 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U575 ( .A(n532), .B(KEYINPUT90), .ZN(G164) );
  NAND2_X1 U576 ( .A1(n526), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U577 ( .A(n520), .B(KEYINPUT67), .ZN(n579) );
  NAND2_X1 U578 ( .A1(G102), .A2(n579), .ZN(n521) );
  XNOR2_X1 U579 ( .A(KEYINPUT89), .B(n521), .ZN(n525) );
  AND2_X1 U580 ( .A1(n571), .A2(G138), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n525), .A2(n524), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G126), .A2(n559), .ZN(n528) );
  NAND2_X1 U583 ( .A1(G114), .A2(n894), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U585 ( .A(KEYINPUT88), .B(n529), .Z(n530) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n652) );
  INV_X1 U587 ( .A(G651), .ZN(n535) );
  NOR2_X1 U588 ( .A1(n652), .A2(n535), .ZN(n664) );
  NAND2_X1 U589 ( .A1(G72), .A2(n664), .ZN(n534) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n666) );
  NAND2_X1 U591 ( .A1(G85), .A2(n666), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n536), .Z(n670) );
  NAND2_X1 U595 ( .A1(G60), .A2(n670), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n652), .A2(G651), .ZN(n537) );
  XNOR2_X1 U597 ( .A(KEYINPUT66), .B(n537), .ZN(n671) );
  NAND2_X1 U598 ( .A1(G47), .A2(n671), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U600 ( .A1(n541), .A2(n540), .ZN(G290) );
  XOR2_X1 U601 ( .A(G2435), .B(G2454), .Z(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT105), .B(G2438), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n543), .B(n542), .ZN(n550) );
  XOR2_X1 U604 ( .A(G2446), .B(G2430), .Z(n545) );
  XNOR2_X1 U605 ( .A(G2451), .B(G2443), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U607 ( .A(n546), .B(G2427), .Z(n548) );
  XNOR2_X1 U608 ( .A(G1348), .B(G1341), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U611 ( .A1(n551), .A2(G14), .ZN(G401) );
  NAND2_X1 U612 ( .A1(G64), .A2(n670), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G52), .A2(n671), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G77), .A2(n664), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G90), .A2(n666), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U619 ( .A1(n558), .A2(n557), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G123), .A2(n559), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n560), .B(KEYINPUT18), .ZN(n569) );
  NAND2_X1 U623 ( .A1(G99), .A2(n561), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G135), .A2(n562), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G111), .A2(n894), .ZN(n565) );
  XNOR2_X1 U627 ( .A(KEYINPUT81), .B(n565), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n937) );
  XNOR2_X1 U630 ( .A(G2096), .B(n937), .ZN(n570) );
  OR2_X1 U631 ( .A1(G2100), .A2(n570), .ZN(G156) );
  INV_X1 U632 ( .A(G120), .ZN(G236) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G113), .A2(n894), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n574), .A2(KEYINPUT69), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G125), .A2(n559), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G101), .A2(n579), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT68), .ZN(n581) );
  XNOR2_X1 U643 ( .A(n581), .B(KEYINPUT23), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U645 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U646 ( .A(G223), .B(KEYINPUT71), .ZN(n845) );
  NAND2_X1 U647 ( .A1(n845), .A2(G567), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U649 ( .A1(n670), .A2(G56), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT14), .B(n586), .Z(n594) );
  XOR2_X1 U651 ( .A(KEYINPUT12), .B(KEYINPUT72), .Z(n588) );
  NAND2_X1 U652 ( .A1(G81), .A2(n666), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n664), .A2(G68), .ZN(n589) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n589), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(KEYINPUT13), .ZN(n593) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(KEYINPUT74), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G43), .A2(n671), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n994) );
  INV_X1 U662 ( .A(n994), .ZN(n598) );
  XOR2_X1 U663 ( .A(G860), .B(KEYINPUT75), .Z(n632) );
  NAND2_X1 U664 ( .A1(n598), .A2(n632), .ZN(G153) );
  NAND2_X1 U665 ( .A1(G79), .A2(n664), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G92), .A2(n666), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U668 ( .A1(G66), .A2(n670), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G54), .A2(n671), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U672 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(n980) );
  INV_X1 U674 ( .A(n980), .ZN(n639) );
  NOR2_X1 U675 ( .A1(G868), .A2(n639), .ZN(n608) );
  INV_X1 U676 ( .A(G868), .ZN(n684) );
  NOR2_X1 U677 ( .A1(G171), .A2(n684), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U679 ( .A(KEYINPUT77), .B(n609), .ZN(G284) );
  NAND2_X1 U680 ( .A1(n666), .A2(G89), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT4), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G76), .A2(n664), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT5), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n670), .A2(G63), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G51), .A2(n671), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT6), .B(n617), .Z(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U692 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U693 ( .A1(G78), .A2(n664), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G91), .A2(n666), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n670), .A2(G65), .ZN(n623) );
  XOR2_X1 U697 ( .A(KEYINPUT70), .B(n623), .Z(n624) );
  NOR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G53), .A2(n671), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(G299) );
  NOR2_X1 U701 ( .A1(G286), .A2(n684), .ZN(n628) );
  XOR2_X1 U702 ( .A(KEYINPUT79), .B(n628), .Z(n630) );
  NOR2_X1 U703 ( .A1(G868), .A2(G299), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(G297) );
  INV_X1 U705 ( .A(G559), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n980), .A2(n633), .ZN(n634) );
  XOR2_X1 U708 ( .A(n634), .B(KEYINPUT16), .Z(n635) );
  XNOR2_X1 U709 ( .A(KEYINPUT80), .B(n635), .ZN(G148) );
  NOR2_X1 U710 ( .A1(G868), .A2(n994), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n639), .A2(G868), .ZN(n636) );
  NOR2_X1 U712 ( .A1(G559), .A2(n636), .ZN(n637) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(G282) );
  NAND2_X1 U714 ( .A1(n639), .A2(G559), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n994), .B(n640), .ZN(n682) );
  NOR2_X1 U716 ( .A1(G860), .A2(n682), .ZN(n648) );
  NAND2_X1 U717 ( .A1(G80), .A2(n664), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G93), .A2(n666), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G67), .A2(n670), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G55), .A2(n671), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  OR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n685) );
  XOR2_X1 U724 ( .A(n685), .B(KEYINPUT82), .Z(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(G145) );
  NAND2_X1 U726 ( .A1(G651), .A2(G74), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G49), .A2(n671), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U729 ( .A1(n670), .A2(n651), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n652), .A2(G87), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(G288) );
  NAND2_X1 U732 ( .A1(n670), .A2(G61), .ZN(n662) );
  NAND2_X1 U733 ( .A1(G86), .A2(n666), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G48), .A2(n671), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n660) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n658) );
  NAND2_X1 U737 ( .A1(n664), .A2(G73), .ZN(n657) );
  XOR2_X1 U738 ( .A(n658), .B(n657), .Z(n659) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U742 ( .A1(G75), .A2(n664), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(KEYINPUT86), .ZN(n669) );
  NAND2_X1 U744 ( .A1(G88), .A2(n666), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT85), .B(n667), .Z(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n675) );
  NAND2_X1 U747 ( .A1(G62), .A2(n670), .ZN(n673) );
  NAND2_X1 U748 ( .A1(G50), .A2(n671), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U750 ( .A1(n675), .A2(n674), .ZN(G166) );
  XOR2_X1 U751 ( .A(n685), .B(G290), .Z(n678) );
  XNOR2_X1 U752 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(G288), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n678), .B(n677), .ZN(n679) );
  INV_X1 U755 ( .A(G299), .ZN(n712) );
  XOR2_X1 U756 ( .A(n679), .B(n712), .Z(n681) );
  XNOR2_X1 U757 ( .A(G305), .B(G166), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n681), .B(n680), .ZN(n873) );
  XNOR2_X1 U759 ( .A(n873), .B(n682), .ZN(n683) );
  NOR2_X1 U760 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U761 ( .A1(G868), .A2(n685), .ZN(n686) );
  NOR2_X1 U762 ( .A1(n687), .A2(n686), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n688) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n688), .Z(n689) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n689), .ZN(n690) );
  XNOR2_X1 U766 ( .A(KEYINPUT21), .B(n690), .ZN(n691) );
  NAND2_X1 U767 ( .A1(n691), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n692) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n692), .Z(n693) );
  NOR2_X1 U771 ( .A1(G218), .A2(n693), .ZN(n694) );
  NAND2_X1 U772 ( .A1(G96), .A2(n694), .ZN(n850) );
  NAND2_X1 U773 ( .A1(n850), .A2(G2106), .ZN(n698) );
  NAND2_X1 U774 ( .A1(G69), .A2(G108), .ZN(n695) );
  NOR2_X1 U775 ( .A1(G236), .A2(n695), .ZN(n696) );
  NAND2_X1 U776 ( .A1(G57), .A2(n696), .ZN(n849) );
  NAND2_X1 U777 ( .A1(n849), .A2(G567), .ZN(n697) );
  NAND2_X1 U778 ( .A1(n698), .A2(n697), .ZN(n927) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n699) );
  NOR2_X1 U780 ( .A1(n927), .A2(n699), .ZN(n848) );
  NAND2_X1 U781 ( .A1(n848), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  NOR2_X1 U783 ( .A1(G1384), .A2(G164), .ZN(n812) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n811) );
  XNOR2_X1 U785 ( .A(n811), .B(KEYINPUT93), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n812), .A2(n700), .ZN(n701) );
  INV_X1 U787 ( .A(n706), .ZN(n702) );
  INV_X2 U788 ( .A(n702), .ZN(n754) );
  NOR2_X1 U789 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U790 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  NOR2_X1 U791 ( .A1(n789), .A2(n704), .ZN(n775) );
  NAND2_X1 U792 ( .A1(n736), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U793 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  INV_X1 U794 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U795 ( .A1(n1008), .A2(n736), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U797 ( .A1(n713), .A2(n712), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(n710), .ZN(n733) );
  NAND2_X1 U799 ( .A1(n713), .A2(n712), .ZN(n731) );
  INV_X1 U800 ( .A(G1341), .ZN(n995) );
  XOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n714) );
  XNOR2_X1 U802 ( .A(KEYINPUT65), .B(n714), .ZN(n719) );
  NAND2_X1 U803 ( .A1(n995), .A2(n719), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n715), .A2(n754), .ZN(n718) );
  INV_X1 U805 ( .A(G1996), .ZN(n956) );
  NOR2_X1 U806 ( .A1(n754), .A2(n956), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n716), .A2(n719), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n726) );
  NOR2_X1 U809 ( .A1(G1996), .A2(n719), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n994), .A2(n720), .ZN(n724) );
  NAND2_X1 U811 ( .A1(G2067), .A2(n736), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n754), .A2(G1348), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n980), .A2(n727), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n729) );
  NOR2_X1 U817 ( .A1(n980), .A2(n727), .ZN(n728) );
  NOR2_X1 U818 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n735) );
  XOR2_X1 U821 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  INV_X1 U822 ( .A(n736), .ZN(n737) );
  NOR2_X1 U823 ( .A1(n961), .A2(n737), .ZN(n739) );
  NOR2_X1 U824 ( .A1(G1961), .A2(n702), .ZN(n738) );
  NOR2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U826 ( .A(KEYINPUT95), .B(n740), .ZN(n746) );
  NAND2_X1 U827 ( .A1(n746), .A2(G171), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n742), .A2(n741), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n754), .A2(G2084), .ZN(n763) );
  NOR2_X1 U830 ( .A1(n766), .A2(n763), .ZN(n743) );
  NAND2_X1 U831 ( .A1(G8), .A2(n743), .ZN(n744) );
  XNOR2_X1 U832 ( .A(KEYINPUT30), .B(n744), .ZN(n745) );
  NOR2_X1 U833 ( .A1(G168), .A2(n745), .ZN(n748) );
  NOR2_X1 U834 ( .A1(G171), .A2(n746), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n752), .A2(n751), .ZN(n764) );
  NAND2_X1 U838 ( .A1(G286), .A2(n764), .ZN(n753) );
  XNOR2_X1 U839 ( .A(n753), .B(KEYINPUT98), .ZN(n760) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n789), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n754), .A2(G2090), .ZN(n755) );
  NOR2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U843 ( .A(KEYINPUT99), .B(n757), .Z(n758) );
  NAND2_X1 U844 ( .A1(n758), .A2(G303), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U847 ( .A(n762), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U848 ( .A1(G8), .A2(n763), .ZN(n768) );
  INV_X1 U849 ( .A(n764), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n770), .A2(n769), .ZN(n778) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U854 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n778), .A2(n772), .ZN(n773) );
  NAND2_X1 U856 ( .A1(n789), .A2(n773), .ZN(n774) );
  NOR2_X1 U857 ( .A1(n775), .A2(n519), .ZN(n794) );
  NAND2_X1 U858 ( .A1(G288), .A2(G1976), .ZN(n776) );
  XOR2_X1 U859 ( .A(KEYINPUT100), .B(n776), .Z(n990) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NOR2_X1 U861 ( .A1(G1971), .A2(G303), .ZN(n777) );
  NOR2_X1 U862 ( .A1(n785), .A2(n777), .ZN(n988) );
  NAND2_X1 U863 ( .A1(n778), .A2(n988), .ZN(n780) );
  NOR2_X1 U864 ( .A1(KEYINPUT101), .A2(n789), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n990), .A2(n781), .ZN(n782) );
  NOR2_X1 U867 ( .A1(KEYINPUT33), .A2(n782), .ZN(n791) );
  INV_X1 U868 ( .A(KEYINPUT101), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n785), .A2(KEYINPUT33), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n785), .A2(KEYINPUT101), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U874 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U875 ( .A1(n792), .A2(n977), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n794), .A2(n793), .ZN(n826) );
  XOR2_X1 U877 ( .A(G1986), .B(G290), .Z(n984) );
  NAND2_X1 U878 ( .A1(G119), .A2(n559), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G95), .A2(n561), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U881 ( .A1(G107), .A2(n894), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G131), .A2(n562), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U884 ( .A1(n800), .A2(n799), .ZN(n906) );
  AND2_X1 U885 ( .A1(n906), .A2(G1991), .ZN(n810) );
  NAND2_X1 U886 ( .A1(G129), .A2(n559), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G117), .A2(n894), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U889 ( .A1(n561), .A2(G105), .ZN(n803) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n803), .Z(n804) );
  NOR2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U892 ( .A(KEYINPUT92), .B(n806), .ZN(n808) );
  NAND2_X1 U893 ( .A1(G141), .A2(n562), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n913) );
  AND2_X1 U895 ( .A1(G1996), .A2(n913), .ZN(n809) );
  NOR2_X1 U896 ( .A1(n810), .A2(n809), .ZN(n828) );
  NAND2_X1 U897 ( .A1(n984), .A2(n828), .ZN(n813) );
  NOR2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n839) );
  NAND2_X1 U899 ( .A1(n813), .A2(n839), .ZN(n824) );
  NAND2_X1 U900 ( .A1(G104), .A2(n561), .ZN(n815) );
  NAND2_X1 U901 ( .A1(G140), .A2(n562), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U903 ( .A(KEYINPUT34), .B(n816), .ZN(n822) );
  NAND2_X1 U904 ( .A1(n559), .A2(G128), .ZN(n817) );
  XOR2_X1 U905 ( .A(KEYINPUT91), .B(n817), .Z(n819) );
  NAND2_X1 U906 ( .A1(n894), .A2(G116), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U908 ( .A(KEYINPUT35), .B(n820), .Z(n821) );
  NOR2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U910 ( .A(KEYINPUT36), .B(n823), .Z(n916) );
  XOR2_X1 U911 ( .A(G2067), .B(KEYINPUT37), .Z(n838) );
  AND2_X1 U912 ( .A1(n916), .A2(n838), .ZN(n934) );
  NAND2_X1 U913 ( .A1(n934), .A2(n839), .ZN(n827) );
  AND2_X1 U914 ( .A1(n824), .A2(n827), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n843) );
  INV_X1 U916 ( .A(n827), .ZN(n837) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n913), .ZN(n946) );
  INV_X1 U918 ( .A(n828), .ZN(n933) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n829) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n906), .ZN(n940) );
  NOR2_X1 U921 ( .A1(n829), .A2(n940), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT103), .B(n830), .Z(n831) );
  NOR2_X1 U923 ( .A1(n933), .A2(n831), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT104), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n946), .A2(n833), .ZN(n834) );
  XNOR2_X1 U926 ( .A(KEYINPUT39), .B(n834), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n835), .A2(n839), .ZN(n836) );
  OR2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n841) );
  NOR2_X1 U929 ( .A1(n916), .A2(n838), .ZN(n936) );
  NAND2_X1 U930 ( .A1(n936), .A2(n839), .ZN(n840) );
  AND2_X1 U931 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U932 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U933 ( .A(n844), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U936 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U938 ( .A1(n848), .A2(n847), .ZN(G188) );
  XOR2_X1 U939 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  XOR2_X1 U940 ( .A(G108), .B(KEYINPUT120), .Z(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  NOR2_X1 U943 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n851), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U945 ( .A(G261), .ZN(G325) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1991), .Z(n853) );
  XNOR2_X1 U947 ( .A(G1981), .B(G1996), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U949 ( .A(n854), .B(KEYINPUT110), .Z(n856) );
  XNOR2_X1 U950 ( .A(G1976), .B(G1971), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U952 ( .A(G1986), .B(G1956), .Z(n858) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1961), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U955 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U956 ( .A(KEYINPUT111), .B(G2474), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n862), .B(n861), .ZN(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(G2678), .Z(n864) );
  XNOR2_X1 U959 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n866) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U964 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(n872) );
  XOR2_X1 U967 ( .A(G2078), .B(G2084), .Z(n871) );
  XNOR2_X1 U968 ( .A(n872), .B(n871), .ZN(G227) );
  XOR2_X1 U969 ( .A(n873), .B(G286), .Z(n875) );
  XNOR2_X1 U970 ( .A(G171), .B(n980), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U972 ( .A(n876), .B(n994), .Z(n877) );
  NOR2_X1 U973 ( .A1(G37), .A2(n877), .ZN(G397) );
  NAND2_X1 U974 ( .A1(n559), .A2(G124), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G100), .A2(n561), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G112), .A2(n894), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G136), .A2(n562), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(G162) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G106), .A2(n561), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G142), .A2(n562), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n893) );
  NAND2_X1 U987 ( .A1(n559), .A2(G130), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n889), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G118), .A2(n894), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n911) );
  NAND2_X1 U992 ( .A1(G127), .A2(n559), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n897), .B(KEYINPUT47), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G139), .A2(n562), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G103), .A2(n561), .ZN(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT115), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n928) );
  XOR2_X1 U1001 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n937), .B(n905), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n906), .B(G162), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n928), .B(n909), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G164), .B(G160), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n917), .B(n916), .Z(n918) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  XNOR2_X1 U1016 ( .A(KEYINPUT118), .B(n920), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n927), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT117), .B(n921), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n922), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n925), .A2(G395), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n926), .B(KEYINPUT119), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(n927), .ZN(G319) );
  INV_X1 U1025 ( .A(G57), .ZN(G237) );
  INV_X1 U1026 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1027 ( .A(G164), .B(G2078), .ZN(n931) );
  XOR2_X1 U1028 ( .A(G2072), .B(n928), .Z(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT121), .B(n929), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT50), .ZN(n944) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n942) );
  XOR2_X1 U1033 ( .A(G2084), .B(G160), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n949) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n947), .Z(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(KEYINPUT122), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n951), .B(KEYINPUT52), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(KEYINPUT55), .A2(n952), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT123), .B(n953), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1048 ( .A(G2067), .B(G26), .Z(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G28), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2072), .B(G33), .Z(n958) );
  XNOR2_X1 U1051 ( .A(n956), .B(G32), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(n961), .B(G27), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G1991), .B(G25), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n966), .B(KEYINPUT53), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G35), .B(G2090), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT55), .B(n972), .ZN(n974) );
  INV_X1 U1065 ( .A(G29), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n975), .A2(G11), .ZN(n1030) );
  INV_X1 U1068 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1069 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n976) );
  XNOR2_X1 U1070 ( .A(n1026), .B(n976), .ZN(n1001) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT57), .ZN(n999) );
  XNOR2_X1 U1074 ( .A(G301), .B(G1961), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n980), .B(G1348), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n993) );
  NAND2_X1 U1077 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G299), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(n991), .Z(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n997) );
  XOR2_X1 U1085 ( .A(n995), .B(n994), .Z(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1028) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n1005) );
  XNOR2_X1 U1090 ( .A(G1976), .B(G23), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1023) );
  XOR2_X1 U1096 ( .A(G1961), .B(G5), .Z(n1018) );
  XNOR2_X1 U1097 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G19), .B(G1341), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT126), .B(G1966), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(G21), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

