

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n518), .B(KEYINPUT23), .ZN(n519) );
  NOR2_X1 U552 ( .A1(n616), .A2(n615), .ZN(n617) );
  INV_X1 U553 ( .A(KEYINPUT100), .ZN(n630) );
  INV_X1 U554 ( .A(KEYINPUT66), .ZN(n518) );
  AND2_X1 U555 ( .A1(n524), .A2(G2104), .ZN(n902) );
  NOR2_X1 U556 ( .A1(G2104), .A2(n524), .ZN(n898) );
  NOR2_X1 U557 ( .A1(G651), .A2(n575), .ZN(n805) );
  XNOR2_X1 U558 ( .A(n520), .B(n519), .ZN(n523) );
  XNOR2_X1 U559 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n761) );
  NOR2_X1 U560 ( .A1(n528), .A2(n527), .ZN(G160) );
  INV_X1 U561 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U562 ( .A1(G101), .A2(n902), .ZN(n520) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n521), .Z(n901) );
  NAND2_X1 U565 ( .A1(G137), .A2(n901), .ZN(n522) );
  NAND2_X1 U566 ( .A1(n523), .A2(n522), .ZN(n528) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U568 ( .A1(G113), .A2(n897), .ZN(n526) );
  NAND2_X1 U569 ( .A1(G125), .A2(n898), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U571 ( .A1(G114), .A2(n897), .ZN(n530) );
  NAND2_X1 U572 ( .A1(G126), .A2(n898), .ZN(n529) );
  AND2_X1 U573 ( .A1(n530), .A2(n529), .ZN(n532) );
  NAND2_X1 U574 ( .A1(G102), .A2(n902), .ZN(n531) );
  AND2_X1 U575 ( .A1(n532), .A2(n531), .ZN(n534) );
  NAND2_X1 U576 ( .A1(n901), .A2(G138), .ZN(n533) );
  AND2_X1 U577 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U578 ( .A(KEYINPUT93), .B(n535), .Z(G164) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n536) );
  XOR2_X1 U580 ( .A(KEYINPUT65), .B(n536), .Z(n802) );
  NAND2_X1 U581 ( .A1(G91), .A2(n802), .ZN(n538) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n575) );
  INV_X1 U583 ( .A(G651), .ZN(n539) );
  NOR2_X1 U584 ( .A1(n575), .A2(n539), .ZN(n809) );
  NAND2_X1 U585 ( .A1(G78), .A2(n809), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n543) );
  NOR2_X1 U587 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n540), .Z(n801) );
  NAND2_X1 U589 ( .A1(G65), .A2(n801), .ZN(n541) );
  XNOR2_X1 U590 ( .A(KEYINPUT69), .B(n541), .ZN(n542) );
  NOR2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U592 ( .A1(n805), .A2(G53), .ZN(n544) );
  NAND2_X1 U593 ( .A1(n545), .A2(n544), .ZN(G299) );
  NAND2_X1 U594 ( .A1(G64), .A2(n801), .ZN(n546) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n546), .Z(n553) );
  NAND2_X1 U596 ( .A1(G90), .A2(n802), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G77), .A2(n809), .ZN(n547) );
  NAND2_X1 U598 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U599 ( .A(n549), .B(KEYINPUT9), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G52), .A2(n805), .ZN(n550) );
  NAND2_X1 U601 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U602 ( .A1(n553), .A2(n552), .ZN(G171) );
  NAND2_X1 U603 ( .A1(n802), .A2(G89), .ZN(n554) );
  XNOR2_X1 U604 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G76), .A2(n809), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U607 ( .A(n557), .B(KEYINPUT5), .ZN(n562) );
  NAND2_X1 U608 ( .A1(G63), .A2(n801), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G51), .A2(n805), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U612 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U613 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U614 ( .A1(G62), .A2(n801), .ZN(n565) );
  NAND2_X1 U615 ( .A1(G88), .A2(n802), .ZN(n564) );
  NAND2_X1 U616 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n809), .A2(G75), .ZN(n566) );
  XOR2_X1 U618 ( .A(KEYINPUT84), .B(n566), .Z(n567) );
  NOR2_X1 U619 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U620 ( .A1(n805), .A2(G50), .ZN(n569) );
  NAND2_X1 U621 ( .A1(n570), .A2(n569), .ZN(G303) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G49), .A2(n805), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U626 ( .A1(n801), .A2(n573), .ZN(n574) );
  XNOR2_X1 U627 ( .A(n574), .B(KEYINPUT80), .ZN(n577) );
  NAND2_X1 U628 ( .A1(G87), .A2(n575), .ZN(n576) );
  NAND2_X1 U629 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U630 ( .A(KEYINPUT81), .B(n578), .Z(G288) );
  NAND2_X1 U631 ( .A1(n809), .A2(G73), .ZN(n580) );
  XNOR2_X1 U632 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n579) );
  XNOR2_X1 U633 ( .A(n580), .B(n579), .ZN(n587) );
  NAND2_X1 U634 ( .A1(G61), .A2(n801), .ZN(n582) );
  NAND2_X1 U635 ( .A1(G86), .A2(n802), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U637 ( .A1(G48), .A2(n805), .ZN(n583) );
  XNOR2_X1 U638 ( .A(KEYINPUT83), .B(n583), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U641 ( .A1(G85), .A2(n802), .ZN(n589) );
  NAND2_X1 U642 ( .A1(G72), .A2(n809), .ZN(n588) );
  NAND2_X1 U643 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U644 ( .A1(G60), .A2(n801), .ZN(n591) );
  NAND2_X1 U645 ( .A1(G47), .A2(n805), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U647 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(n594), .ZN(G290) );
  XOR2_X1 U649 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n667) );
  NAND2_X1 U650 ( .A1(G54), .A2(n805), .ZN(n601) );
  NAND2_X1 U651 ( .A1(G92), .A2(n802), .ZN(n596) );
  NAND2_X1 U652 ( .A1(G79), .A2(n809), .ZN(n595) );
  NAND2_X1 U653 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U654 ( .A1(n801), .A2(G66), .ZN(n597) );
  XOR2_X1 U655 ( .A(KEYINPUT74), .B(n597), .Z(n598) );
  NOR2_X1 U656 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U657 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U658 ( .A(n602), .B(KEYINPUT15), .ZN(n985) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n709) );
  INV_X1 U660 ( .A(n709), .ZN(n603) );
  NOR2_X2 U661 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NAND2_X2 U662 ( .A1(n603), .A2(n708), .ZN(n656) );
  INV_X1 U663 ( .A(G1996), .ZN(n953) );
  NOR2_X1 U664 ( .A1(n656), .A2(n953), .ZN(n604) );
  XNOR2_X1 U665 ( .A(n604), .B(KEYINPUT26), .ZN(n616) );
  NAND2_X1 U666 ( .A1(G56), .A2(n801), .ZN(n605) );
  XOR2_X1 U667 ( .A(KEYINPUT14), .B(n605), .Z(n611) );
  NAND2_X1 U668 ( .A1(n802), .A2(G81), .ZN(n606) );
  XNOR2_X1 U669 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U670 ( .A1(G68), .A2(n809), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U672 ( .A(KEYINPUT13), .B(n609), .Z(n610) );
  NOR2_X1 U673 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U674 ( .A1(n805), .A2(G43), .ZN(n612) );
  NAND2_X1 U675 ( .A1(n613), .A2(n612), .ZN(n978) );
  AND2_X1 U676 ( .A1(n656), .A2(G1341), .ZN(n614) );
  OR2_X1 U677 ( .A1(n978), .A2(n614), .ZN(n615) );
  XNOR2_X1 U678 ( .A(KEYINPUT64), .B(n617), .ZN(n629) );
  NAND2_X1 U679 ( .A1(n985), .A2(n629), .ZN(n621) );
  INV_X1 U680 ( .A(n656), .ZN(n641) );
  NOR2_X1 U681 ( .A1(n641), .A2(G1348), .ZN(n619) );
  NOR2_X1 U682 ( .A1(G2067), .A2(n656), .ZN(n618) );
  NOR2_X1 U683 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U684 ( .A1(n621), .A2(n620), .ZN(n628) );
  INV_X1 U685 ( .A(G299), .ZN(n975) );
  INV_X1 U686 ( .A(G2072), .ZN(n622) );
  OR2_X1 U687 ( .A1(n656), .A2(n622), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n623), .B(KEYINPUT27), .ZN(n626) );
  NAND2_X1 U689 ( .A1(G1956), .A2(n656), .ZN(n624) );
  XNOR2_X1 U690 ( .A(KEYINPUT99), .B(n624), .ZN(n625) );
  NOR2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n634) );
  NOR2_X1 U692 ( .A1(n975), .A2(n634), .ZN(n627) );
  XOR2_X1 U693 ( .A(n627), .B(KEYINPUT28), .Z(n636) );
  AND2_X1 U694 ( .A1(n628), .A2(n636), .ZN(n633) );
  NOR2_X1 U695 ( .A1(n985), .A2(n629), .ZN(n631) );
  XNOR2_X1 U696 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n638) );
  AND2_X1 U698 ( .A1(n975), .A2(n634), .ZN(n635) );
  NAND2_X1 U699 ( .A1(n636), .A2(n635), .ZN(n637) );
  AND2_X1 U700 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U701 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n639) );
  XNOR2_X1 U702 ( .A(n640), .B(n639), .ZN(n645) );
  XNOR2_X1 U703 ( .A(KEYINPUT25), .B(G2078), .ZN(n955) );
  NOR2_X1 U704 ( .A1(n656), .A2(n955), .ZN(n643) );
  INV_X1 U705 ( .A(G1961), .ZN(n1001) );
  NOR2_X1 U706 ( .A1(n641), .A2(n1001), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U708 ( .A1(n646), .A2(G171), .ZN(n644) );
  NAND2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n670) );
  NOR2_X1 U710 ( .A1(G171), .A2(n646), .ZN(n654) );
  INV_X1 U711 ( .A(G8), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n647), .A2(G1966), .ZN(n648) );
  AND2_X1 U713 ( .A1(n656), .A2(n648), .ZN(n672) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n656), .ZN(n668) );
  NOR2_X1 U715 ( .A1(n672), .A2(n668), .ZN(n649) );
  XNOR2_X1 U716 ( .A(KEYINPUT102), .B(n649), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n650), .A2(G8), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U719 ( .A1(G168), .A2(n652), .ZN(n653) );
  NOR2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT31), .B(n655), .Z(n669) );
  NAND2_X1 U722 ( .A1(G8), .A2(n656), .ZN(n703) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n703), .ZN(n658) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n656), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(G303), .ZN(n661) );
  AND2_X1 U727 ( .A1(n669), .A2(n661), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n670), .A2(n660), .ZN(n664) );
  INV_X1 U729 ( .A(n661), .ZN(n662) );
  OR2_X1 U730 ( .A1(n662), .A2(G286), .ZN(n663) );
  AND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(n676) );
  NAND2_X1 U734 ( .A1(G8), .A2(n668), .ZN(n674) );
  AND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n701) );
  NOR2_X1 U739 ( .A1(G288), .A2(G1976), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT104), .ZN(n681) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n681), .A2(n678), .ZN(n989) );
  NAND2_X1 U743 ( .A1(n701), .A2(n989), .ZN(n680) );
  INV_X1 U744 ( .A(KEYINPUT105), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n680), .B(n679), .ZN(n691) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U747 ( .A(KEYINPUT33), .ZN(n693) );
  INV_X1 U748 ( .A(n703), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n693), .A2(n683), .ZN(n684) );
  XOR2_X1 U751 ( .A(n684), .B(KEYINPUT106), .Z(n692) );
  AND2_X1 U752 ( .A1(n980), .A2(n692), .ZN(n688) );
  NOR2_X1 U753 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XOR2_X1 U754 ( .A(n685), .B(KEYINPUT24), .Z(n686) );
  OR2_X1 U755 ( .A1(n703), .A2(n686), .ZN(n695) );
  XNOR2_X1 U756 ( .A(G1981), .B(G305), .ZN(n995) );
  AND2_X1 U757 ( .A1(n695), .A2(n995), .ZN(n698) );
  INV_X1 U758 ( .A(n698), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U760 ( .A1(n703), .A2(n689), .ZN(n690) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n707) );
  INV_X1 U762 ( .A(n692), .ZN(n694) );
  OR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n696) );
  AND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n705) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n742) );
  NOR2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U773 ( .A(n710), .B(KEYINPUT94), .ZN(n757) );
  XOR2_X1 U774 ( .A(G1986), .B(G290), .Z(n984) );
  XOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .Z(n711) );
  XOR2_X1 U776 ( .A(KEYINPUT95), .B(n711), .Z(n746) );
  XNOR2_X1 U777 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G140), .A2(n901), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G104), .A2(n902), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U781 ( .A(n715), .B(n714), .ZN(n720) );
  NAND2_X1 U782 ( .A1(G116), .A2(n897), .ZN(n717) );
  NAND2_X1 U783 ( .A1(G128), .A2(n898), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U785 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U787 ( .A(KEYINPUT36), .B(n721), .Z(n889) );
  AND2_X1 U788 ( .A1(n746), .A2(n889), .ZN(n753) );
  NAND2_X1 U789 ( .A1(G141), .A2(n901), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G117), .A2(n897), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U792 ( .A1(n902), .A2(G105), .ZN(n724) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U795 ( .A1(n898), .A2(G129), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n908) );
  NAND2_X1 U797 ( .A1(G1996), .A2(n908), .ZN(n729) );
  XNOR2_X1 U798 ( .A(n729), .B(KEYINPUT98), .ZN(n738) );
  NAND2_X1 U799 ( .A1(G131), .A2(n901), .ZN(n731) );
  NAND2_X1 U800 ( .A1(G107), .A2(n897), .ZN(n730) );
  NAND2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U802 ( .A1(G95), .A2(n902), .ZN(n732) );
  XNOR2_X1 U803 ( .A(KEYINPUT97), .B(n732), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U805 ( .A1(n898), .A2(G119), .ZN(n735) );
  NAND2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n894) );
  NAND2_X1 U807 ( .A1(G1991), .A2(n894), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n749) );
  NOR2_X1 U809 ( .A1(n753), .A2(n749), .ZN(n928) );
  NAND2_X1 U810 ( .A1(n984), .A2(n928), .ZN(n745) );
  NAND2_X1 U811 ( .A1(n757), .A2(n745), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n742), .A2(n739), .ZN(n741) );
  INV_X1 U813 ( .A(KEYINPUT107), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n742), .A2(KEYINPUT107), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n760) );
  NAND2_X1 U817 ( .A1(n745), .A2(KEYINPUT107), .ZN(n756) );
  NOR2_X1 U818 ( .A1(n746), .A2(n889), .ZN(n946) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n908), .ZN(n933) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U821 ( .A1(G1991), .A2(n894), .ZN(n926) );
  NOR2_X1 U822 ( .A1(n747), .A2(n926), .ZN(n748) );
  NOR2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n933), .A2(n750), .ZN(n751) );
  XOR2_X1 U825 ( .A(KEYINPUT39), .B(n751), .Z(n752) );
  NOR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n946), .A2(n754), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U831 ( .A(n762), .B(n761), .ZN(G329) );
  XNOR2_X1 U832 ( .A(G2454), .B(G2427), .ZN(n772) );
  XOR2_X1 U833 ( .A(KEYINPUT110), .B(G2430), .Z(n764) );
  XNOR2_X1 U834 ( .A(G2443), .B(G2451), .ZN(n763) );
  XNOR2_X1 U835 ( .A(n764), .B(n763), .ZN(n768) );
  XOR2_X1 U836 ( .A(G2446), .B(KEYINPUT109), .Z(n766) );
  XNOR2_X1 U837 ( .A(G1348), .B(G1341), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U839 ( .A(n768), .B(n767), .Z(n770) );
  XNOR2_X1 U840 ( .A(G2435), .B(G2438), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U842 ( .A(n772), .B(n771), .ZN(n773) );
  AND2_X1 U843 ( .A1(n773), .A2(G14), .ZN(G401) );
  AND2_X1 U844 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U845 ( .A(G57), .ZN(G237) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U848 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U849 ( .A(G223), .B(KEYINPUT71), .ZN(n844) );
  NAND2_X1 U850 ( .A1(n844), .A2(G567), .ZN(n775) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n781) );
  OR2_X1 U853 ( .A1(n978), .A2(n781), .ZN(n776) );
  XNOR2_X1 U854 ( .A(KEYINPUT72), .B(n776), .ZN(G153) );
  XNOR2_X1 U855 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n778) );
  OR2_X1 U857 ( .A1(n985), .A2(G868), .ZN(n777) );
  NAND2_X1 U858 ( .A1(n778), .A2(n777), .ZN(G284) );
  INV_X1 U859 ( .A(G868), .ZN(n824) );
  NOR2_X1 U860 ( .A1(G286), .A2(n824), .ZN(n780) );
  NOR2_X1 U861 ( .A1(G868), .A2(G299), .ZN(n779) );
  NOR2_X1 U862 ( .A1(n780), .A2(n779), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n781), .A2(G559), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n782), .A2(n985), .ZN(n783) );
  XNOR2_X1 U865 ( .A(n783), .B(KEYINPUT75), .ZN(n784) );
  XOR2_X1 U866 ( .A(KEYINPUT16), .B(n784), .Z(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n978), .ZN(n785) );
  XNOR2_X1 U868 ( .A(KEYINPUT76), .B(n785), .ZN(n788) );
  NAND2_X1 U869 ( .A1(G868), .A2(n985), .ZN(n786) );
  NOR2_X1 U870 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U871 ( .A1(n788), .A2(n787), .ZN(G282) );
  NAND2_X1 U872 ( .A1(G99), .A2(n902), .ZN(n795) );
  NAND2_X1 U873 ( .A1(G135), .A2(n901), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G111), .A2(n897), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n898), .A2(G123), .ZN(n791) );
  XOR2_X1 U877 ( .A(KEYINPUT18), .B(n791), .Z(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT77), .ZN(n930) );
  XNOR2_X1 U881 ( .A(G2096), .B(n930), .ZN(n798) );
  INV_X1 U882 ( .A(G2100), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(G156) );
  NAND2_X1 U884 ( .A1(G559), .A2(n985), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(n978), .ZN(n822) );
  XNOR2_X1 U886 ( .A(KEYINPUT78), .B(n822), .ZN(n800) );
  NOR2_X1 U887 ( .A1(G860), .A2(n800), .ZN(n812) );
  NAND2_X1 U888 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G55), .A2(n805), .ZN(n806) );
  XNOR2_X1 U892 ( .A(KEYINPUT79), .B(n806), .ZN(n807) );
  NOR2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n809), .A2(G80), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n825) );
  XOR2_X1 U896 ( .A(n812), .B(n825), .Z(G145) );
  INV_X1 U897 ( .A(G303), .ZN(G166) );
  XOR2_X1 U898 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n814) );
  XNOR2_X1 U899 ( .A(G166), .B(KEYINPUT19), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U901 ( .A(KEYINPUT88), .B(n815), .ZN(n817) );
  XNOR2_X1 U902 ( .A(G288), .B(KEYINPUT85), .ZN(n816) );
  XNOR2_X1 U903 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U904 ( .A(n818), .B(G290), .ZN(n819) );
  XNOR2_X1 U905 ( .A(n819), .B(G305), .ZN(n820) );
  XNOR2_X1 U906 ( .A(n975), .B(n820), .ZN(n821) );
  XNOR2_X1 U907 ( .A(n821), .B(n825), .ZN(n914) );
  XNOR2_X1 U908 ( .A(n822), .B(n914), .ZN(n823) );
  NAND2_X1 U909 ( .A1(n823), .A2(G868), .ZN(n827) );
  NAND2_X1 U910 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U911 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(n828), .Z(n829) );
  NAND2_X1 U914 ( .A1(G2090), .A2(n829), .ZN(n830) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n830), .ZN(n831) );
  NAND2_X1 U916 ( .A1(n831), .A2(G2072), .ZN(G158) );
  XOR2_X1 U917 ( .A(KEYINPUT89), .B(G44), .Z(n832) );
  XNOR2_X1 U918 ( .A(KEYINPUT3), .B(n832), .ZN(G218) );
  XOR2_X1 U919 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U920 ( .A1(G219), .A2(G220), .ZN(n834) );
  XNOR2_X1 U921 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n833) );
  XNOR2_X1 U922 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U923 ( .A(KEYINPUT22), .B(n835), .ZN(n836) );
  NOR2_X1 U924 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U925 ( .A1(G96), .A2(n837), .ZN(n849) );
  NAND2_X1 U926 ( .A1(n849), .A2(G2106), .ZN(n842) );
  NAND2_X1 U927 ( .A1(G69), .A2(G120), .ZN(n838) );
  NOR2_X1 U928 ( .A1(G237), .A2(n838), .ZN(n839) );
  NAND2_X1 U929 ( .A1(G108), .A2(n839), .ZN(n848) );
  NAND2_X1 U930 ( .A1(G567), .A2(n848), .ZN(n840) );
  XNOR2_X1 U931 ( .A(KEYINPUT92), .B(n840), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n842), .A2(n841), .ZN(n850) );
  NAND2_X1 U933 ( .A1(G483), .A2(G661), .ZN(n843) );
  NOR2_X1 U934 ( .A1(n850), .A2(n843), .ZN(n847) );
  NAND2_X1 U935 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(G188) );
  XNOR2_X1 U941 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  INV_X1 U947 ( .A(n850), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2474), .B(G1976), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1956), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(KEYINPUT113), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1991), .B(G1996), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G1981), .B(G1971), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G229) );
  XOR2_X1 U960 ( .A(G2096), .B(KEYINPUT112), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2090), .B(KEYINPUT43), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n864), .B(KEYINPUT42), .Z(n866) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2072), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(G2678), .B(G2100), .Z(n868) );
  XNOR2_X1 U967 ( .A(G2078), .B(G2084), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(G227) );
  NAND2_X1 U970 ( .A1(G124), .A2(n898), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT44), .B(n871), .Z(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT115), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G112), .A2(n897), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G136), .A2(n901), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G100), .A2(n902), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n880) );
  XNOR2_X1 U980 ( .A(KEYINPUT118), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n893) );
  NAND2_X1 U982 ( .A1(G139), .A2(n901), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G103), .A2(n902), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n897), .A2(G115), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT117), .B(n883), .Z(n885) );
  NAND2_X1 U987 ( .A1(n898), .A2(G127), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n939) );
  XOR2_X1 U991 ( .A(G162), .B(n939), .Z(n891) );
  XNOR2_X1 U992 ( .A(G164), .B(n889), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n894), .B(n930), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n912) );
  NAND2_X1 U997 ( .A1(G118), .A2(n897), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n901), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n902), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n905), .B(KEYINPUT45), .Z(n906) );
  NOR2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(G160), .B(n910), .Z(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G286), .B(n978), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1011 ( .A(G171), .B(n985), .Z(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n920), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT119), .B(n922), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n931), .Z(n936) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1032 ( .A(KEYINPUT121), .B(n937), .Z(n944) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT122), .B(n938), .ZN(n941) );
  XOR2_X1 U1035 ( .A(G2072), .B(n939), .Z(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT50), .B(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n971), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n949), .A2(G29), .ZN(n1029) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n962) );
  XOR2_X1 U1048 ( .A(G1991), .B(G25), .Z(n952) );
  NAND2_X1 U1049 ( .A1(n952), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n953), .B(G32), .ZN(n957) );
  XOR2_X1 U1051 ( .A(G27), .B(KEYINPUT123), .Z(n954) );
  XNOR2_X1 U1052 ( .A(n955), .B(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT124), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT125), .B(n963), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT53), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1060 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n971), .B(n970), .ZN(n973) );
  INV_X1 U1064 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n974), .ZN(n1027) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1068 ( .A(n975), .B(G1956), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1071 ( .A(G1341), .B(n978), .Z(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n992) );
  XNOR2_X1 U1075 ( .A(G171), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n985), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT127), .B(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n998) );
  XOR2_X1 U1081 ( .A(G1966), .B(G168), .Z(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n993), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT57), .B(n996), .Z(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1025) );
  INV_X1 U1087 ( .A(G16), .ZN(n1023) );
  XNOR2_X1 U1088 ( .A(G5), .B(n1001), .ZN(n1018) );
  XOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G4), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G20), .B(G1956), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1009), .B(KEYINPUT60), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(G1986), .B(G24), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(G1976), .B(G23), .Z(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

