//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT73), .B(G902), .Z(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G953), .A3(new_n187), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT21), .B(G898), .Z(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G214), .B1(G237), .B2(G902), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(KEYINPUT68), .A3(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT5), .ZN(new_n206));
  AOI211_X1 g020(.A(new_n206), .B(new_n197), .C1(new_n200), .C2(new_n201), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n197), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G113), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n205), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT77), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  OAI21_X1  g033(.A(G107), .B1(new_n212), .B2(KEYINPUT3), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(KEYINPUT77), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n212), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(G104), .B2(new_n216), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n224), .A3(new_n226), .A4(new_n212), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G101), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n211), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G110), .B(G122), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT83), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT8), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n232), .B(KEYINPUT83), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n230), .A2(new_n222), .ZN(new_n240));
  INV_X1    g054(.A(new_n208), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n202), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n208), .B2(new_n197), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n242), .A2(new_n244), .B1(new_n202), .B2(new_n204), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n231), .A2(new_n239), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n240), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT77), .B(G107), .ZN(new_n252));
  OR2_X1    g066(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n220), .B(new_n221), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n254), .A2(G101), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(G101), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n254), .B2(G101), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n202), .B2(new_n204), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n196), .A2(KEYINPUT68), .A3(G119), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT68), .B1(new_n196), .B2(G119), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n262), .A2(new_n263), .B1(new_n196), .B2(G119), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n203), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n260), .A3(new_n203), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n251), .B(new_n234), .C1(new_n259), .C2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n231), .A2(new_n239), .A3(new_n246), .A4(KEYINPUT88), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n249), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n188), .A2(G224), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT87), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n274));
  INV_X1    g088(.A(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G146), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n276), .A2(new_n278), .A3(new_n279), .A4(KEYINPUT65), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT0), .ZN(new_n285));
  INV_X1    g099(.A(G128), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n279), .B1(new_n276), .B2(new_n278), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n282), .A2(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G125), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n277), .B(G146), .C1(new_n286), .C2(KEYINPUT1), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(new_n275), .A3(G143), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n302));
  XNOR2_X1  g116(.A(G143), .B(G146), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n286), .A2(KEYINPUT1), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND4_X1   g119(.A1(new_n302), .A2(new_n304), .A3(new_n276), .A4(new_n278), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n299), .B(new_n301), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT86), .B1(new_n307), .B2(G125), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n296), .A2(new_n300), .A3(new_n297), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n300), .B1(new_n296), .B2(new_n297), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n276), .A3(new_n278), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT66), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n303), .A2(new_n302), .A3(new_n304), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n315), .A3(new_n316), .A4(new_n292), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n274), .B1(new_n295), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n271), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n295), .A2(KEYINPUT7), .A3(new_n273), .A4(new_n318), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n273), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n293), .B(KEYINPUT85), .ZN(new_n324));
  INV_X1    g138(.A(new_n318), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n295), .A2(new_n273), .A3(new_n318), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n259), .A2(new_n268), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n242), .A2(new_n244), .ZN(new_n330));
  AND4_X1   g144(.A1(new_n205), .A2(new_n330), .A3(new_n222), .A4(new_n230), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n236), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n269), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n334));
  INV_X1    g148(.A(new_n268), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n258), .A2(new_n257), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n254), .A2(G101), .A3(new_n255), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n234), .B1(new_n339), .B2(new_n251), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT6), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n334), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n331), .B1(new_n335), .B2(new_n338), .ZN(new_n343));
  NOR4_X1   g157(.A1(new_n343), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n234), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n328), .B(new_n333), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n322), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT89), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n322), .A2(new_n345), .A3(new_n349), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n195), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G469), .ZN(new_n354));
  INV_X1    g168(.A(new_n190), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  INV_X1    g170(.A(G227), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G953), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n356), .B(new_n358), .Z(new_n359));
  AOI21_X1  g173(.A(new_n298), .B1(new_n313), .B2(new_n314), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT80), .B1(new_n240), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n296), .B(new_n297), .C1(new_n305), .C2(new_n306), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n222), .A4(new_n230), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n250), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n290), .A2(new_n289), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT65), .B1(new_n303), .B2(new_n279), .ZN(new_n371));
  INV_X1    g185(.A(new_n283), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n259), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n376), .A3(new_n366), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(G137), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(G137), .ZN(new_n382));
  INV_X1    g196(.A(G137), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT11), .A3(G134), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  INV_X1    g200(.A(G131), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n384), .A3(new_n387), .A4(new_n382), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n386), .A2(new_n388), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n368), .A2(new_n391), .A3(new_n375), .A4(new_n377), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n359), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n240), .A2(new_n315), .A3(new_n311), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n365), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n389), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT12), .ZN(new_n399));
  AND4_X1   g213(.A1(new_n392), .A2(new_n359), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n354), .B(new_n355), .C1(new_n393), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G902), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n354), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n359), .B(KEYINPUT76), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n376), .B1(new_n365), .B2(new_n366), .ZN(new_n406));
  AOI211_X1 g220(.A(KEYINPUT81), .B(KEYINPUT10), .C1(new_n361), .C2(new_n364), .ZN(new_n407));
  NOR4_X1   g221(.A1(new_n406), .A2(new_n407), .A3(new_n389), .A4(new_n374), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n397), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n390), .A2(new_n392), .A3(new_n359), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G469), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n404), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT9), .B(G234), .Z(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n188), .A3(G214), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n277), .ZN(new_n419));
  NOR2_X1   g233(.A1(G237), .A2(G953), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(G143), .A3(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n387), .A3(new_n421), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT91), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n292), .A2(KEYINPUT16), .A3(G140), .ZN(new_n428));
  XNOR2_X1  g242(.A(G125), .B(G140), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G146), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n430), .A2(G146), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n423), .A2(new_n436), .A3(new_n424), .A4(new_n425), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n427), .A2(new_n434), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n429), .B(new_n275), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n387), .ZN(new_n441));
  OAI221_X1 g255(.A(new_n439), .B1(new_n422), .B2(new_n441), .C1(new_n423), .C2(new_n440), .ZN(new_n442));
  XOR2_X1   g256(.A(G113), .B(G122), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT90), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(G104), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n438), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n438), .B2(new_n442), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n402), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT94), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT93), .B(G475), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(new_n402), .C1(new_n446), .C2(new_n447), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n445), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n429), .B(KEYINPUT19), .Z(new_n455));
  OAI21_X1  g269(.A(new_n431), .B1(new_n455), .B2(G146), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n423), .A2(new_n425), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n442), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n438), .A2(new_n442), .A3(new_n445), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(KEYINPUT92), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n462), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n453), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(G116), .B(G122), .Z(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(new_n252), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n196), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  OAI211_X1 g287(.A(G107), .B(new_n473), .C1(new_n471), .C2(KEYINPUT14), .ZN(new_n474));
  XNOR2_X1  g288(.A(G128), .B(G143), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT95), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n476), .A2(new_n380), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n380), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n472), .B(new_n474), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n380), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n471), .B(new_n252), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(KEYINPUT13), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n277), .A2(G128), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(G134), .C1(KEYINPUT13), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G217), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n415), .A2(new_n486), .A3(G953), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n479), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n479), .B2(new_n485), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT96), .B(new_n355), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n490), .B(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n470), .A2(new_n493), .ZN(new_n494));
  AND4_X1   g308(.A1(new_n353), .A2(new_n413), .A3(new_n416), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n199), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n286), .A2(G119), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G110), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G110), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n199), .A2(KEYINPUT23), .A3(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n502), .A2(new_n503), .B1(new_n199), .B2(G128), .ZN(new_n504));
  OAI221_X1 g318(.A(new_n500), .B1(new_n501), .B2(new_n504), .C1(new_n432), .C2(new_n433), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(new_n501), .B1(new_n498), .B2(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n429), .A2(new_n275), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n431), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT22), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G137), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n505), .B(new_n514), .C1(new_n509), .C2(new_n510), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n355), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT25), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n486), .B1(new_n355), .B2(G234), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n516), .A2(new_n521), .A3(new_n355), .A4(new_n517), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n520), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  INV_X1    g344(.A(new_n382), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n380), .A2(G137), .ZN(new_n532));
  OAI21_X1  g346(.A(G131), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n388), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n307), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n291), .A2(new_n389), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n268), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT70), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n307), .A2(new_n535), .B1(new_n291), .B2(new_n389), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n268), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n536), .A2(new_n544), .A3(new_n537), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n536), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n335), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(G101), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n420), .A2(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n543), .A2(new_n547), .A3(new_n554), .A4(new_n551), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n530), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT28), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n538), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n540), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n335), .ZN(new_n561));
  AND4_X1   g375(.A1(new_n541), .A2(new_n268), .A3(new_n536), .A4(new_n537), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n541), .B1(new_n540), .B2(new_n268), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n564), .B2(KEYINPUT28), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n551), .B(KEYINPUT72), .Z(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI22_X1  g381(.A1(new_n565), .A2(new_n567), .B1(KEYINPUT31), .B2(new_n552), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n529), .B(new_n402), .C1(new_n556), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT32), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n391), .A2(new_n373), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n534), .B1(new_n311), .B2(new_n315), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT30), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n536), .A2(new_n544), .A3(new_n537), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n335), .A2(new_n575), .B1(new_n539), .B2(new_n542), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n554), .B1(new_n576), .B2(new_n551), .ZN(new_n577));
  AND4_X1   g391(.A1(new_n554), .A2(new_n543), .A3(new_n547), .A4(new_n551), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT31), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n539), .A2(new_n542), .B1(new_n560), .B2(new_n335), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n558), .B1(new_n580), .B2(new_n557), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n562), .A2(new_n563), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n268), .B1(new_n573), .B2(new_n574), .ZN(new_n583));
  INV_X1    g397(.A(new_n551), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n581), .A2(new_n566), .B1(new_n585), .B2(new_n530), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n529), .A4(new_n402), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n576), .B2(new_n551), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n551), .B(new_n558), .C1(new_n580), .C2(new_n557), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n566), .A2(KEYINPUT29), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n565), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n190), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n591), .B1(new_n598), .B2(new_n529), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n593), .A2(new_n594), .B1(new_n565), .B2(new_n596), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT74), .B(G472), .C1(new_n600), .C2(new_n190), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n528), .B1(new_n590), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n495), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n413), .A2(new_n416), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n190), .B1(new_n579), .B2(new_n586), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n527), .B(new_n569), .C1(new_n609), .C2(new_n529), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n612), .A2(KEYINPUT98), .A3(new_n416), .A4(new_n413), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n346), .A2(new_n347), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n322), .A2(new_n345), .A3(new_n348), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n194), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n488), .A2(new_n489), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n491), .A3(new_n355), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n479), .A2(new_n485), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n620), .A2(KEYINPUT33), .A3(new_n625), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n355), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n623), .B1(new_n629), .B2(G478), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n470), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n615), .A2(KEYINPUT99), .A3(new_n194), .A4(new_n616), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n619), .A2(new_n633), .A3(new_n193), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n614), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AND2_X1   g452(.A1(new_n453), .A2(new_n469), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n466), .A2(new_n462), .A3(new_n468), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n464), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n639), .A2(new_n493), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n619), .A2(new_n193), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n614), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n511), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n525), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n523), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n569), .B(new_n650), .C1(new_n609), .C2(new_n529), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n495), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AOI22_X1  g469(.A1(new_n570), .A2(new_n589), .B1(new_n599), .B2(new_n601), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n608), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n619), .A2(new_n634), .A3(new_n650), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n189), .B(KEYINPUT101), .Z(new_n660));
  INV_X1    g474(.A(new_n191), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  INV_X1    g481(.A(new_n416), .ZN(new_n668));
  INV_X1    g482(.A(new_n359), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n406), .A2(new_n407), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n391), .B1(new_n670), .B2(new_n375), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n671), .B2(new_n408), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n392), .A2(new_n359), .A3(new_n397), .A4(new_n399), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n190), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n403), .B1(new_n674), .B2(new_n354), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n668), .B1(new_n675), .B2(new_n412), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n663), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT106), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n351), .A2(new_n352), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT102), .Z(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n493), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n632), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n523), .A3(new_n649), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n553), .A2(new_n555), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n566), .A2(new_n564), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n529), .B1(new_n690), .B2(KEYINPUT103), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n689), .B(new_n691), .C1(KEYINPUT103), .C2(new_n690), .ZN(new_n692));
  NAND2_X1  g506(.A1(G472), .A2(G902), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n688), .B1(new_n696), .B2(new_n590), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n684), .A2(new_n194), .A3(new_n685), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT38), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n683), .B(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n194), .A4(new_n697), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n679), .A2(new_n680), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n681), .A2(new_n699), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NAND3_X1  g520(.A1(new_n630), .A2(new_n470), .A3(new_n664), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n659), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  OAI21_X1  g524(.A(new_n355), .B1(new_n393), .B2(new_n400), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n416), .A3(new_n401), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n656), .A2(new_n528), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n635), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  INV_X1    g532(.A(new_n643), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND2_X1  g535(.A1(new_n672), .A2(new_n673), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n354), .B1(new_n722), .B2(new_n355), .ZN(new_n723));
  AOI211_X1 g537(.A(G469), .B(new_n190), .C1(new_n672), .C2(new_n673), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n619), .A3(new_n416), .A4(new_n634), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n656), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n494), .A2(new_n193), .A3(new_n650), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NAND4_X1  g545(.A1(new_n619), .A2(new_n193), .A3(new_n634), .A4(new_n687), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n713), .A2(new_n610), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NAND2_X1  g550(.A1(new_n652), .A2(new_n708), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n726), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n619), .A2(new_n634), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n723), .A2(new_n724), .A3(new_n668), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n651), .A2(new_n707), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  INV_X1    g559(.A(new_n194), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n682), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n411), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n411), .A2(new_n748), .ZN(new_n750));
  OAI211_X1 g564(.A(G469), .B(new_n410), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n668), .B1(new_n751), .B2(new_n675), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n603), .A2(new_n708), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT110), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n603), .A2(new_n665), .A3(new_n747), .A4(new_n752), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  OAI211_X1 g576(.A(KEYINPUT45), .B(new_n410), .C1(new_n749), .C2(new_n750), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n410), .B2(new_n411), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n354), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n404), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n401), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  INV_X1    g584(.A(new_n766), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n403), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n773), .A3(new_n401), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n632), .A2(new_n630), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT43), .Z(new_n777));
  OAI21_X1  g591(.A(new_n569), .B1(new_n609), .B2(new_n529), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(KEYINPUT44), .A3(new_n778), .A4(new_n650), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n416), .A3(new_n677), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n778), .A3(new_n650), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n747), .B1(new_n782), .B2(KEYINPUT44), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n383), .ZN(G39));
  XNOR2_X1  g599(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n775), .B2(new_n416), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n775), .A2(new_n416), .A3(new_n786), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n708), .A3(new_n747), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n590), .A2(new_n602), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n527), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(G140), .Z(G42));
  INV_X1    g609(.A(new_n701), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n696), .A2(new_n527), .A3(new_n590), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n776), .A2(new_n746), .A3(new_n668), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n725), .B(KEYINPUT49), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n791), .A2(new_n741), .A3(new_n527), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n741), .A2(new_n612), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n802), .A2(new_n635), .B1(new_n803), .B2(new_n732), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n727), .A2(new_n729), .B1(new_n714), .B2(new_n719), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n756), .A2(new_n757), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n470), .A2(new_n686), .A3(KEYINPUT113), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT113), .B1(new_n470), .B2(new_n686), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n808), .B(new_n809), .C1(new_n632), .C2(new_n631), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n611), .A2(new_n613), .A3(new_n353), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n495), .B1(new_n603), .B2(new_n652), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n639), .A2(new_n641), .A3(new_n650), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n814), .A2(new_n682), .A3(new_n746), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n493), .A2(new_n663), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n791), .A2(new_n676), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n752), .A2(new_n742), .A3(new_n747), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n761), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n697), .A2(new_n739), .A3(new_n664), .A4(new_n752), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n657), .B(new_n658), .C1(new_n665), .C2(new_n708), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n744), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n744), .A2(new_n822), .A3(KEYINPUT52), .A4(new_n823), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n827), .A2(KEYINPUT114), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n801), .A2(new_n821), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(KEYINPUT53), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n832), .B2(new_n801), .ZN(new_n836));
  AOI211_X1 g650(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n821), .C2(new_n831), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n813), .A2(new_n819), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n807), .B1(KEYINPUT116), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n801), .B1(new_n820), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n829), .A3(new_n828), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n777), .A2(new_n660), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n610), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n739), .A3(new_n741), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n188), .A2(G952), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n741), .A2(new_n747), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n189), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n797), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n633), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n846), .A2(new_n850), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n528), .A3(new_n656), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  AOI211_X1 g670(.A(new_n849), .B(new_n853), .C1(new_n856), .C2(KEYINPUT48), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n834), .A2(new_n845), .A3(new_n848), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n725), .A2(new_n668), .ZN(new_n859));
  INV_X1    g673(.A(new_n789), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n787), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n747), .A3(new_n847), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n852), .A2(new_n632), .A3(new_n631), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n701), .A2(new_n846), .A3(new_n194), .A4(new_n803), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT50), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n854), .A2(new_n651), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT51), .Z(new_n868));
  NOR3_X1   g682(.A1(new_n855), .A2(KEYINPUT117), .A3(KEYINPUT48), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n858), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(G952), .A2(G953), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n800), .B1(new_n870), .B2(new_n871), .ZN(G75));
  NAND4_X1  g686(.A1(new_n791), .A2(new_n741), .A3(new_n619), .A4(new_n634), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n873), .A2(new_n728), .B1(new_n802), .B2(new_n643), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n804), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n840), .A2(new_n756), .A3(new_n875), .A4(new_n757), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n827), .B2(new_n826), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT115), .B1(new_n877), .B2(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n832), .A2(new_n835), .A3(new_n801), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n844), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n190), .A3(new_n348), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n333), .B1(new_n342), .B2(new_n344), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT118), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n328), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n188), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n887), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n882), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n888), .A2(new_n895), .A3(new_n890), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n403), .B(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n839), .B1(new_n838), .B2(new_n844), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n839), .A2(new_n878), .A3(new_n844), .A4(new_n879), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT120), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n722), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n355), .B1(new_n838), .B2(new_n844), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n771), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n889), .B1(new_n905), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n466), .A2(new_n468), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n889), .ZN(G60));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT59), .Z(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n834), .B2(new_n845), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n627), .B2(new_n628), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n899), .A2(new_n900), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n627), .A2(new_n628), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n915), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n917), .A2(new_n920), .A3(new_n889), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT60), .Z(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n838), .B2(new_n844), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n889), .B1(new_n925), .B2(new_n648), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n524), .B2(new_n925), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n926), .B(KEYINPUT61), .C1(new_n524), .C2(new_n925), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(G66));
  NAND2_X1  g745(.A1(new_n192), .A2(G224), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G953), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n813), .A2(new_n874), .A3(new_n804), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT122), .Z(new_n936));
  INV_X1    g750(.A(G898), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n885), .B1(new_n937), .B2(G953), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n936), .B(new_n938), .ZN(G69));
  XOR2_X1   g753(.A(new_n575), .B(new_n455), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n357), .B2(new_n662), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n744), .A2(new_n823), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n705), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g760(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n678), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n603), .A3(new_n747), .A4(new_n810), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n950), .C1(new_n793), .C2(new_n790), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n705), .A2(new_n945), .A3(new_n953), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n951), .A2(new_n784), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n943), .B1(new_n955), .B2(new_n188), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n739), .A2(new_n603), .A3(new_n687), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n775), .A2(new_n416), .A3(new_n677), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n758), .A2(new_n958), .A3(new_n761), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n790), .B2(new_n793), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n784), .B2(new_n944), .ZN(new_n964));
  OAI211_X1 g778(.A(KEYINPUT124), .B(new_n945), .C1(new_n780), .C2(new_n783), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT126), .B(G900), .ZN(new_n971));
  OAI22_X1  g785(.A1(new_n970), .A2(G953), .B1(new_n942), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n956), .B1(new_n972), .B2(new_n940), .ZN(G72));
  INV_X1    g787(.A(new_n576), .ZN(new_n974));
  INV_X1    g788(.A(new_n934), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n951), .A2(new_n784), .A3(new_n975), .A4(new_n954), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n693), .B(KEYINPUT63), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n974), .B(new_n551), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(new_n584), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n689), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n889), .B1(new_n833), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n966), .A2(new_n934), .A3(new_n969), .ZN(new_n983));
  INV_X1    g797(.A(new_n977), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n983), .A2(KEYINPUT127), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT127), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n974), .A2(new_n551), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n987), .B2(new_n988), .ZN(G57));
endmodule


