

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786;

  NAND2_X1 U373 ( .A1(n639), .A2(n776), .ZN(n756) );
  NOR2_X1 U374 ( .A1(n603), .A2(n633), .ZN(n605) );
  AND2_X1 U375 ( .A1(n644), .A2(n756), .ZN(n680) );
  INV_X1 U376 ( .A(n680), .ZN(n693) );
  BUF_X1 U377 ( .A(n483), .Z(n775) );
  NOR2_X1 U378 ( .A1(n481), .A2(n482), .ZN(n566) );
  NOR2_X2 U379 ( .A1(n578), .A2(n784), .ZN(n579) );
  INV_X1 U380 ( .A(n724), .ZN(n367) );
  XNOR2_X2 U381 ( .A(n519), .B(n430), .ZN(n671) );
  NOR2_X1 U382 ( .A1(n601), .A2(n600), .ZN(n410) );
  NOR2_X2 U383 ( .A1(n553), .A2(n723), .ZN(n622) );
  INV_X1 U384 ( .A(n626), .ZN(n734) );
  AND2_X1 U385 ( .A1(n408), .A2(n638), .ZN(n407) );
  NOR2_X1 U386 ( .A1(n783), .A2(n612), .ZN(n613) );
  NOR2_X1 U387 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U388 ( .A(n410), .B(n357), .ZN(n427) );
  NOR2_X1 U389 ( .A1(n581), .A2(n711), .ZN(n531) );
  XNOR2_X1 U390 ( .A(n593), .B(n356), .ZN(n601) );
  AND2_X1 U391 ( .A1(n580), .A2(n711), .ZN(n746) );
  NOR2_X1 U392 ( .A1(n744), .A2(n745), .ZN(n533) );
  XNOR2_X1 U393 ( .A(n557), .B(n556), .ZN(n707) );
  XNOR2_X1 U394 ( .A(n500), .B(n499), .ZN(n549) );
  NAND2_X1 U395 ( .A1(n400), .A2(n397), .ZN(n364) );
  XNOR2_X1 U396 ( .A(n470), .B(n440), .ZN(n695) );
  XNOR2_X1 U397 ( .A(n426), .B(n443), .ZN(n640) );
  XNOR2_X1 U398 ( .A(G125), .B(G146), .ZN(n488) );
  XNOR2_X2 U399 ( .A(n458), .B(n457), .ZN(n596) );
  NAND2_X1 U400 ( .A1(n640), .A2(KEYINPUT84), .ZN(n380) );
  NAND2_X1 U401 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U402 ( .A1(n723), .A2(KEYINPUT108), .ZN(n366) );
  AND2_X1 U403 ( .A1(n370), .A2(n369), .ZN(n368) );
  OR2_X1 U404 ( .A1(n695), .A2(n398), .ZN(n397) );
  NAND2_X1 U405 ( .A1(n442), .A2(n399), .ZN(n398) );
  AND2_X1 U406 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U407 ( .A1(n403), .A2(G902), .ZN(n401) );
  INV_X1 U408 ( .A(KEYINPUT47), .ZN(n417) );
  NOR2_X1 U409 ( .A1(n746), .A2(n417), .ZN(n412) );
  AND2_X1 U410 ( .A1(n632), .A2(n631), .ZN(n637) );
  INV_X1 U411 ( .A(G237), .ZN(n472) );
  NAND2_X1 U412 ( .A1(n379), .A2(n378), .ZN(n377) );
  AND2_X1 U413 ( .A1(n381), .A2(n380), .ZN(n378) );
  NAND2_X1 U414 ( .A1(n641), .A2(n382), .ZN(n381) );
  XNOR2_X1 U415 ( .A(n488), .B(n446), .ZN(n507) );
  XOR2_X1 U416 ( .A(KEYINPUT10), .B(G140), .Z(n446) );
  XNOR2_X1 U417 ( .A(n470), .B(n469), .ZN(n663) );
  XOR2_X1 U418 ( .A(n507), .B(n447), .Z(n669) );
  XNOR2_X1 U419 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U420 ( .A(G128), .B(G110), .ZN(n453) );
  XNOR2_X1 U421 ( .A(G122), .B(G107), .ZN(n495) );
  XNOR2_X1 U422 ( .A(n707), .B(n558), .ZN(n580) );
  XNOR2_X1 U423 ( .A(n529), .B(n686), .ZN(n555) );
  NAND2_X1 U424 ( .A1(n364), .A2(KEYINPUT1), .ZN(n372) );
  NAND2_X1 U425 ( .A1(n383), .A2(n359), .ZN(n394) );
  OR2_X1 U426 ( .A1(n659), .A2(G210), .ZN(n395) );
  AND2_X1 U427 ( .A1(n386), .A2(n391), .ZN(n385) );
  NAND2_X1 U428 ( .A1(n693), .A2(n393), .ZN(n386) );
  AND2_X1 U429 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U430 ( .A1(G953), .A2(G237), .ZN(n503) );
  XNOR2_X1 U431 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n487) );
  XNOR2_X1 U432 ( .A(G902), .B(KEYINPUT91), .ZN(n426) );
  XNOR2_X1 U433 ( .A(n579), .B(KEYINPUT86), .ZN(n421) );
  XNOR2_X1 U434 ( .A(n361), .B(n358), .ZN(n578) );
  XNOR2_X1 U435 ( .A(G131), .B(G143), .ZN(n508) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n475) );
  INV_X1 U437 ( .A(KEYINPUT45), .ZN(n428) );
  XNOR2_X1 U438 ( .A(n425), .B(n445), .ZN(n728) );
  AND2_X1 U439 ( .A1(n455), .A2(G221), .ZN(n425) );
  AND2_X1 U440 ( .A1(n421), .A2(n582), .ZN(n757) );
  INV_X1 U441 ( .A(G146), .ZN(n439) );
  XNOR2_X1 U442 ( .A(G107), .B(G140), .ZN(n433) );
  AND2_X1 U443 ( .A1(n659), .A2(G210), .ZN(n396) );
  INV_X1 U444 ( .A(KEYINPUT89), .ZN(n550) );
  XNOR2_X1 U445 ( .A(n611), .B(KEYINPUT35), .ZN(n616) );
  INV_X1 U446 ( .A(KEYINPUT34), .ZN(n607) );
  AND2_X1 U447 ( .A1(n362), .A2(n644), .ZN(n665) );
  XNOR2_X1 U448 ( .A(n454), .B(n450), .ZN(n423) );
  XNOR2_X1 U449 ( .A(n528), .B(n527), .ZN(n688) );
  NAND2_X1 U450 ( .A1(n525), .A2(n524), .ZN(n528) );
  AND2_X1 U451 ( .A1(n363), .A2(n644), .ZN(n649) );
  XNOR2_X1 U452 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n628) );
  NOR2_X1 U453 ( .A1(n563), .A2(n555), .ZN(n557) );
  XNOR2_X1 U454 ( .A(n409), .B(KEYINPUT107), .ZN(n654) );
  NOR2_X1 U455 ( .A1(n601), .A2(n595), .ZN(n409) );
  NAND2_X1 U456 ( .A1(n429), .A2(n635), .ZN(n700) );
  INV_X1 U457 ( .A(n601), .ZN(n429) );
  AND2_X1 U458 ( .A1(n392), .A2(n389), .ZN(n388) );
  NAND2_X1 U459 ( .A1(n372), .A2(n371), .ZN(n724) );
  NOR2_X1 U460 ( .A1(n626), .A2(n625), .ZN(n352) );
  XOR2_X1 U461 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n353) );
  INV_X1 U462 ( .A(n723), .ZN(n374) );
  AND2_X1 U463 ( .A1(n397), .A2(n373), .ZN(n354) );
  INV_X1 U464 ( .A(G902), .ZN(n399) );
  AND2_X1 U465 ( .A1(n582), .A2(KEYINPUT2), .ZN(n355) );
  XOR2_X1 U466 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n356) );
  INV_X1 U467 ( .A(KEYINPUT1), .ZN(n373) );
  XOR2_X1 U468 ( .A(n602), .B(KEYINPUT32), .Z(n357) );
  INV_X1 U469 ( .A(n659), .ZN(n393) );
  XOR2_X1 U470 ( .A(n570), .B(KEYINPUT70), .Z(n358) );
  INV_X1 U471 ( .A(KEYINPUT84), .ZN(n382) );
  AND2_X1 U472 ( .A1(n395), .A2(n684), .ZN(n359) );
  AND2_X1 U473 ( .A1(n380), .A2(n382), .ZN(n360) );
  NAND2_X1 U474 ( .A1(n569), .A2(n568), .ZN(n361) );
  AND2_X1 U475 ( .A1(n756), .A2(G472), .ZN(n362) );
  AND2_X1 U476 ( .A1(n756), .A2(G475), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n695), .A2(n403), .ZN(n402) );
  XNOR2_X2 U478 ( .A(n671), .B(n439), .ZN(n470) );
  NAND2_X1 U479 ( .A1(n367), .A2(n374), .ZN(n625) );
  NAND2_X1 U480 ( .A1(n368), .A2(n365), .ZN(n603) );
  NAND2_X1 U481 ( .A1(n723), .A2(KEYINPUT108), .ZN(n369) );
  NAND2_X1 U482 ( .A1(n724), .A2(KEYINPUT108), .ZN(n370) );
  NAND2_X1 U483 ( .A1(n400), .A2(n397), .ZN(n553) );
  NAND2_X1 U484 ( .A1(n354), .A2(n400), .ZN(n371) );
  NAND2_X1 U485 ( .A1(n375), .A2(n757), .ZN(n643) );
  NAND2_X1 U486 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U487 ( .A1(n759), .A2(n360), .ZN(n376) );
  INV_X1 U488 ( .A(n759), .ZN(n379) );
  XNOR2_X2 U489 ( .A(n404), .B(n428), .ZN(n759) );
  NAND2_X1 U490 ( .A1(n680), .A2(n396), .ZN(n383) );
  NAND2_X1 U491 ( .A1(n388), .A2(n384), .ZN(G51) );
  NAND2_X1 U492 ( .A1(n387), .A2(n385), .ZN(n384) );
  INV_X1 U493 ( .A(n394), .ZN(n387) );
  NAND2_X1 U494 ( .A1(n693), .A2(n390), .ZN(n389) );
  NOR2_X1 U495 ( .A1(n659), .A2(n391), .ZN(n390) );
  INV_X1 U496 ( .A(n661), .ZN(n391) );
  NAND2_X1 U497 ( .A1(n394), .A2(n661), .ZN(n392) );
  INV_X1 U498 ( .A(n442), .ZN(n403) );
  NAND2_X1 U499 ( .A1(n407), .A2(n405), .ZN(n404) );
  NAND2_X1 U500 ( .A1(n406), .A2(n615), .ZN(n405) );
  NAND2_X1 U501 ( .A1(n613), .A2(n614), .ZN(n406) );
  NAND2_X1 U502 ( .A1(n620), .A2(n621), .ZN(n408) );
  NAND2_X1 U503 ( .A1(n427), .A2(n654), .ZN(n619) );
  NAND2_X1 U504 ( .A1(n414), .A2(n411), .ZN(n419) );
  NAND2_X1 U505 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U506 ( .A(n712), .ZN(n413) );
  NAND2_X1 U507 ( .A1(n746), .A2(n417), .ZN(n415) );
  NAND2_X1 U508 ( .A1(n712), .A2(n417), .ZN(n416) );
  XNOR2_X1 U509 ( .A(n418), .B(KEYINPUT77), .ZN(n567) );
  NAND2_X1 U510 ( .A1(n419), .A2(n710), .ZN(n418) );
  NAND2_X1 U511 ( .A1(n421), .A2(n355), .ZN(n420) );
  XNOR2_X1 U512 ( .A(n420), .B(KEYINPUT85), .ZN(n639) );
  NOR2_X1 U513 ( .A1(n681), .A2(G902), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n669), .B(n422), .ZN(n681) );
  XNOR2_X1 U515 ( .A(n451), .B(n423), .ZN(n422) );
  NAND2_X1 U516 ( .A1(n424), .A2(n534), .ZN(n535) );
  INV_X1 U517 ( .A(n728), .ZN(n424) );
  XNOR2_X1 U518 ( .A(n427), .B(G119), .ZN(G21) );
  INV_X2 U519 ( .A(G953), .ZN(n483) );
  XNOR2_X1 U520 ( .A(n519), .B(n521), .ZN(n523) );
  BUF_X2 U521 ( .A(n549), .Z(n574) );
  XNOR2_X2 U522 ( .A(n574), .B(KEYINPUT38), .ZN(n742) );
  XNOR2_X2 U523 ( .A(n560), .B(KEYINPUT19), .ZN(n590) );
  XOR2_X1 U524 ( .A(G131), .B(KEYINPUT4), .Z(n430) );
  INV_X1 U525 ( .A(n746), .ZN(n631) );
  INV_X1 U526 ( .A(KEYINPUT48), .ZN(n570) );
  XNOR2_X1 U527 ( .A(n520), .B(n353), .ZN(n521) );
  INV_X1 U528 ( .A(G134), .ZN(n438) );
  INV_X1 U529 ( .A(KEYINPUT24), .ZN(n452) );
  XNOR2_X1 U530 ( .A(n441), .B(n692), .ZN(n442) );
  INV_X1 U531 ( .A(KEYINPUT105), .ZN(n558) );
  INV_X1 U532 ( .A(KEYINPUT104), .ZN(n556) );
  XNOR2_X1 U533 ( .A(n629), .B(n628), .ZN(n718) );
  INV_X1 U534 ( .A(KEYINPUT60), .ZN(n652) );
  XNOR2_X1 U535 ( .A(n653), .B(n652), .ZN(G60) );
  XNOR2_X1 U536 ( .A(KEYINPUT80), .B(G110), .ZN(n431) );
  XNOR2_X1 U537 ( .A(n431), .B(G104), .ZN(n770) );
  XNOR2_X1 U538 ( .A(KEYINPUT67), .B(G101), .ZN(n461) );
  XNOR2_X1 U539 ( .A(n770), .B(n461), .ZN(n491) );
  XOR2_X1 U540 ( .A(G137), .B(KEYINPUT69), .Z(n447) );
  INV_X1 U541 ( .A(n447), .ZN(n435) );
  NAND2_X1 U542 ( .A1(n483), .A2(G227), .ZN(n432) );
  XOR2_X1 U543 ( .A(n433), .B(n432), .Z(n434) );
  XNOR2_X1 U544 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U545 ( .A(n491), .B(n436), .ZN(n440) );
  INV_X2 U546 ( .A(G143), .ZN(n437) );
  XNOR2_X2 U547 ( .A(n437), .B(G128), .ZN(n485) );
  XNOR2_X2 U548 ( .A(n485), .B(n438), .ZN(n519) );
  XNOR2_X1 U549 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n441) );
  INV_X1 U550 ( .A(G469), .ZN(n692) );
  INV_X1 U551 ( .A(KEYINPUT15), .ZN(n443) );
  NAND2_X1 U552 ( .A1(n640), .A2(G234), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n444), .B(KEYINPUT20), .ZN(n455) );
  INV_X1 U554 ( .A(KEYINPUT21), .ZN(n445) );
  NAND2_X1 U555 ( .A1(n775), .A2(G234), .ZN(n449) );
  XOR2_X1 U556 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n448) );
  XNOR2_X1 U557 ( .A(n449), .B(n448), .ZN(n526) );
  NAND2_X1 U558 ( .A1(G221), .A2(n526), .ZN(n451) );
  XOR2_X1 U559 ( .A(G119), .B(KEYINPUT23), .Z(n450) );
  AND2_X1 U560 ( .A1(G217), .A2(n455), .ZN(n456) );
  XNOR2_X1 U561 ( .A(KEYINPUT25), .B(n456), .ZN(n457) );
  OR2_X2 U562 ( .A1(n728), .A2(n596), .ZN(n723) );
  XNOR2_X1 U563 ( .A(KEYINPUT111), .B(n622), .ZN(n482) );
  XOR2_X1 U564 ( .A(KEYINPUT5), .B(KEYINPUT79), .Z(n460) );
  XNOR2_X1 U565 ( .A(KEYINPUT94), .B(KEYINPUT78), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U567 ( .A(n462), .B(n461), .ZN(n468) );
  NAND2_X1 U568 ( .A1(n503), .A2(G210), .ZN(n464) );
  XNOR2_X1 U569 ( .A(G116), .B(G137), .ZN(n463) );
  XNOR2_X1 U570 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U571 ( .A(KEYINPUT3), .B(G119), .ZN(n465) );
  XNOR2_X1 U572 ( .A(n465), .B(G113), .ZN(n494) );
  XNOR2_X1 U573 ( .A(n466), .B(n494), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U575 ( .A1(n663), .A2(n399), .ZN(n471) );
  INV_X1 U576 ( .A(G472), .ZN(n662) );
  XNOR2_X2 U577 ( .A(n471), .B(n662), .ZN(n626) );
  NAND2_X1 U578 ( .A1(n399), .A2(n472), .ZN(n498) );
  NAND2_X1 U579 ( .A1(n498), .A2(G214), .ZN(n741) );
  NAND2_X1 U580 ( .A1(n734), .A2(n741), .ZN(n473) );
  XNOR2_X1 U581 ( .A(KEYINPUT30), .B(n473), .ZN(n474) );
  INV_X1 U582 ( .A(n474), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n475), .B(KEYINPUT14), .ZN(n477) );
  NAND2_X1 U584 ( .A1(G952), .A2(n477), .ZN(n476) );
  XOR2_X1 U585 ( .A(KEYINPUT92), .B(n476), .Z(n754) );
  NAND2_X1 U586 ( .A1(n754), .A2(n775), .ZN(n587) );
  NAND2_X1 U587 ( .A1(G902), .A2(n477), .ZN(n583) );
  NOR2_X1 U588 ( .A1(G900), .A2(n583), .ZN(n478) );
  NAND2_X1 U589 ( .A1(G953), .A2(n478), .ZN(n479) );
  NAND2_X1 U590 ( .A1(n587), .A2(n479), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n480), .A2(n534), .ZN(n481) );
  NAND2_X1 U592 ( .A1(n483), .A2(G224), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n484), .B(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U594 ( .A(n485), .B(n486), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n492) );
  XNOR2_X1 U597 ( .A(n492), .B(n491), .ZN(n497) );
  XNOR2_X1 U598 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n494), .B(n493), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n495), .B(G116), .ZN(n522) );
  XNOR2_X1 U601 ( .A(n496), .B(n522), .ZN(n772) );
  XNOR2_X1 U602 ( .A(n497), .B(n772), .ZN(n658) );
  INV_X1 U603 ( .A(n640), .ZN(n641) );
  OR2_X2 U604 ( .A1(n658), .A2(n641), .ZN(n500) );
  NAND2_X1 U605 ( .A1(n498), .A2(G210), .ZN(n499) );
  NAND2_X1 U606 ( .A1(n566), .A2(n742), .ZN(n502) );
  INV_X1 U607 ( .A(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U608 ( .A(n502), .B(n501), .ZN(n581) );
  XOR2_X1 U609 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n505) );
  NAND2_X1 U610 ( .A1(G214), .A2(n503), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n507), .B(n506), .ZN(n515) );
  XOR2_X1 U613 ( .A(G104), .B(G113), .Z(n509) );
  XNOR2_X1 U614 ( .A(n509), .B(n508), .ZN(n513) );
  XOR2_X1 U615 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n511) );
  XNOR2_X1 U616 ( .A(G122), .B(KEYINPUT99), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U618 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U619 ( .A(n515), .B(n514), .ZN(n647) );
  NOR2_X1 U620 ( .A1(G902), .A2(n647), .ZN(n517) );
  XNOR2_X1 U621 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n516) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U623 ( .A(G475), .ZN(n645) );
  XNOR2_X1 U624 ( .A(n518), .B(n645), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n520) );
  OR2_X1 U626 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U627 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U628 ( .A1(n526), .A2(G217), .ZN(n527) );
  NAND2_X1 U629 ( .A1(n688), .A2(n399), .ZN(n529) );
  INV_X1 U630 ( .A(G478), .ZN(n686) );
  NAND2_X1 U631 ( .A1(n563), .A2(n555), .ZN(n711) );
  INV_X1 U632 ( .A(KEYINPUT40), .ZN(n530) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n786) );
  INV_X1 U634 ( .A(n555), .ZN(n564) );
  OR2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n744) );
  NAND2_X1 U636 ( .A1(n742), .A2(n741), .ZN(n745) );
  XNOR2_X1 U637 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n763) );
  XNOR2_X1 U639 ( .A(n535), .B(KEYINPUT71), .ZN(n536) );
  NAND2_X1 U640 ( .A1(n596), .A2(n536), .ZN(n545) );
  NOR2_X1 U641 ( .A1(n545), .A2(n626), .ZN(n537) );
  XNOR2_X1 U642 ( .A(n537), .B(KEYINPUT28), .ZN(n539) );
  INV_X1 U643 ( .A(n553), .ZN(n538) );
  NAND2_X1 U644 ( .A1(n539), .A2(n538), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n763), .A2(n559), .ZN(n540) );
  XOR2_X1 U646 ( .A(KEYINPUT42), .B(n540), .Z(n785) );
  NAND2_X1 U647 ( .A1(n786), .A2(n785), .ZN(n543) );
  XOR2_X1 U648 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n541) );
  XNOR2_X1 U649 ( .A(KEYINPUT88), .B(n541), .ZN(n542) );
  XNOR2_X1 U650 ( .A(n543), .B(n542), .ZN(n569) );
  INV_X1 U651 ( .A(KEYINPUT6), .ZN(n544) );
  XNOR2_X1 U652 ( .A(n626), .B(n544), .ZN(n633) );
  NOR2_X1 U653 ( .A1(n633), .A2(n545), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n546), .B(KEYINPUT109), .ZN(n547) );
  NOR2_X1 U655 ( .A1(n711), .A2(n547), .ZN(n571) );
  INV_X1 U656 ( .A(n741), .ZN(n548) );
  NOR2_X2 U657 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X2 U658 ( .A(n551), .B(n550), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n571), .A2(n560), .ZN(n552) );
  XOR2_X1 U660 ( .A(KEYINPUT36), .B(n552), .Z(n554) );
  NAND2_X1 U661 ( .A1(n554), .A2(n367), .ZN(n721) );
  INV_X1 U662 ( .A(n559), .ZN(n562) );
  INV_X1 U663 ( .A(n590), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n562), .A2(n561), .ZN(n712) );
  NAND2_X1 U665 ( .A1(n564), .A2(n563), .ZN(n609) );
  NOR2_X1 U666 ( .A1(n609), .A2(n574), .ZN(n565) );
  NAND2_X1 U667 ( .A1(n566), .A2(n565), .ZN(n710) );
  AND2_X1 U668 ( .A1(n721), .A2(n567), .ZN(n568) );
  NAND2_X1 U669 ( .A1(n571), .A2(n741), .ZN(n572) );
  NOR2_X1 U670 ( .A1(n367), .A2(n572), .ZN(n573) );
  XNOR2_X1 U671 ( .A(n573), .B(KEYINPUT43), .ZN(n576) );
  INV_X1 U672 ( .A(n574), .ZN(n575) );
  NOR2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U674 ( .A(n577), .B(KEYINPUT110), .ZN(n784) );
  OR2_X1 U675 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U676 ( .A(n582), .ZN(n722) );
  INV_X1 U677 ( .A(n583), .ZN(n585) );
  INV_X1 U678 ( .A(G898), .ZN(n584) );
  AND2_X1 U679 ( .A1(n584), .A2(G953), .ZN(n773) );
  NAND2_X1 U680 ( .A1(n585), .A2(n773), .ZN(n586) );
  NAND2_X1 U681 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U682 ( .A(n588), .B(KEYINPUT93), .ZN(n589) );
  NOR2_X2 U683 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X2 U684 ( .A(n591), .B(KEYINPUT0), .ZN(n627) );
  NOR2_X1 U685 ( .A1(n744), .A2(n728), .ZN(n592) );
  NAND2_X1 U686 ( .A1(n627), .A2(n592), .ZN(n593) );
  AND2_X1 U687 ( .A1(n626), .A2(n596), .ZN(n594) );
  NAND2_X1 U688 ( .A1(n724), .A2(n594), .ZN(n595) );
  XNOR2_X1 U689 ( .A(n596), .B(KEYINPUT106), .ZN(n727) );
  INV_X1 U690 ( .A(n727), .ZN(n597) );
  NOR2_X1 U691 ( .A1(n724), .A2(n597), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n598), .A2(n633), .ZN(n599) );
  XNOR2_X1 U693 ( .A(n599), .B(KEYINPUT82), .ZN(n600) );
  INV_X1 U694 ( .A(KEYINPUT81), .ZN(n602) );
  INV_X1 U695 ( .A(KEYINPUT65), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n619), .A2(n617), .ZN(n614) );
  XNOR2_X1 U697 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n604) );
  XNOR2_X1 U698 ( .A(n605), .B(n604), .ZN(n740) );
  INV_X1 U699 ( .A(n627), .ZN(n606) );
  NOR2_X1 U700 ( .A1(n740), .A2(n606), .ZN(n608) );
  XNOR2_X1 U701 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U702 ( .A(n616), .ZN(n783) );
  INV_X1 U703 ( .A(KEYINPUT44), .ZN(n612) );
  OR2_X1 U704 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n615) );
  NAND2_X1 U705 ( .A1(n616), .A2(n612), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n618), .A2(n617), .ZN(n621) );
  INV_X1 U707 ( .A(n619), .ZN(n620) );
  AND2_X1 U708 ( .A1(n622), .A2(n626), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n627), .A2(n623), .ZN(n624) );
  XNOR2_X1 U710 ( .A(KEYINPUT95), .B(n624), .ZN(n703) );
  NAND2_X1 U711 ( .A1(n627), .A2(n352), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n703), .A2(n718), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n630), .B(KEYINPUT97), .ZN(n632) );
  NOR2_X1 U714 ( .A1(n367), .A2(n727), .ZN(n634) );
  AND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n635) );
  INV_X1 U716 ( .A(n700), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  INV_X1 U718 ( .A(n759), .ZN(n776) );
  NAND2_X1 U719 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U721 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U724 ( .A(G952), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n650), .A2(G953), .ZN(n684) );
  NAND2_X1 U726 ( .A1(n651), .A2(n684), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(G110), .ZN(G12) );
  XOR2_X1 U728 ( .A(KEYINPUT83), .B(KEYINPUT90), .Z(n656) );
  XNOR2_X1 U729 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U732 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT87), .ZN(n661) );
  XOR2_X1 U734 ( .A(KEYINPUT62), .B(n663), .Z(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(n684), .ZN(n668) );
  XOR2_X1 U737 ( .A(KEYINPUT113), .B(KEYINPUT63), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G57) );
  XOR2_X1 U739 ( .A(n669), .B(KEYINPUT125), .Z(n670) );
  XOR2_X1 U740 ( .A(n671), .B(n670), .Z(n673) );
  XNOR2_X1 U741 ( .A(n757), .B(n673), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(n775), .ZN(n679) );
  XOR2_X1 U743 ( .A(G227), .B(n673), .Z(n674) );
  NAND2_X1 U744 ( .A1(n674), .A2(G900), .ZN(n675) );
  XOR2_X1 U745 ( .A(KEYINPUT126), .B(n675), .Z(n676) );
  NOR2_X1 U746 ( .A1(n676), .A2(n775), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT127), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(G72) );
  NAND2_X1 U749 ( .A1(n680), .A2(G217), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n681), .B(KEYINPUT124), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n685) );
  INV_X1 U752 ( .A(n684), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n685), .A2(n698), .ZN(G66) );
  NOR2_X1 U754 ( .A1(n693), .A2(n686), .ZN(n690) );
  XOR2_X1 U755 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n687) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n691), .A2(n698), .ZN(G63) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n697) );
  XNOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(G54) );
  XNOR2_X1 U764 ( .A(G101), .B(KEYINPUT114), .ZN(n701) );
  XNOR2_X1 U765 ( .A(n701), .B(n700), .ZN(G3) );
  INV_X1 U766 ( .A(n711), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n703), .A2(n715), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n702), .B(G104), .ZN(G6) );
  XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n705) );
  INV_X1 U770 ( .A(n707), .ZN(n717) );
  NAND2_X1 U771 ( .A1(n703), .A2(n717), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U773 ( .A(G107), .B(n706), .ZN(G9) );
  NOR2_X1 U774 ( .A1(n712), .A2(n707), .ZN(n709) );
  XNOR2_X1 U775 ( .A(G128), .B(KEYINPUT29), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n709), .B(n708), .ZN(G30) );
  XNOR2_X1 U777 ( .A(G143), .B(n710), .ZN(G45) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U779 ( .A(G146), .B(KEYINPUT115), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n714), .B(n713), .ZN(G48) );
  NAND2_X1 U781 ( .A1(n718), .A2(n715), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(G113), .ZN(G15) );
  NAND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U784 ( .A(n719), .B(G116), .ZN(G18) );
  XOR2_X1 U785 ( .A(G125), .B(KEYINPUT37), .Z(n720) );
  XNOR2_X1 U786 ( .A(n721), .B(n720), .ZN(G27) );
  XOR2_X1 U787 ( .A(G134), .B(n722), .Z(G36) );
  XOR2_X1 U788 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n726) );
  NAND2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U790 ( .A(n726), .B(n725), .ZN(n732) );
  XOR2_X1 U791 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n730) );
  NAND2_X1 U792 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U793 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U794 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U795 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U796 ( .A1(n352), .A2(n735), .ZN(n736) );
  XOR2_X1 U797 ( .A(n736), .B(KEYINPUT51), .Z(n737) );
  XNOR2_X1 U798 ( .A(KEYINPUT118), .B(n737), .ZN(n738) );
  NOR2_X1 U799 ( .A1(n763), .A2(n738), .ZN(n739) );
  XOR2_X1 U800 ( .A(KEYINPUT119), .B(n739), .Z(n751) );
  NOR2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n744), .A2(n743), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U804 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U805 ( .A1(n740), .A2(n749), .ZN(n750) );
  NOR2_X1 U806 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U807 ( .A(KEYINPUT52), .B(n752), .Z(n753) );
  NAND2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT120), .ZN(n767) );
  INV_X1 U810 ( .A(n756), .ZN(n762) );
  INV_X1 U811 ( .A(n757), .ZN(n758) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U813 ( .A1(n760), .A2(KEYINPUT2), .ZN(n761) );
  NOR2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n765) );
  NOR2_X1 U815 ( .A1(n740), .A2(n763), .ZN(n764) );
  NOR2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U817 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U818 ( .A1(n768), .A2(G953), .ZN(n769) );
  XNOR2_X1 U819 ( .A(n769), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U820 ( .A(n770), .B(G101), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(n774) );
  NOR2_X1 U822 ( .A1(n774), .A2(n773), .ZN(n782) );
  NAND2_X1 U823 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U824 ( .A1(G953), .A2(G224), .ZN(n777) );
  XNOR2_X1 U825 ( .A(KEYINPUT61), .B(n777), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(G898), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U828 ( .A(n782), .B(n781), .ZN(G69) );
  XOR2_X1 U829 ( .A(G122), .B(n783), .Z(G24) );
  XOR2_X1 U830 ( .A(G140), .B(n784), .Z(G42) );
  XNOR2_X1 U831 ( .A(G137), .B(n785), .ZN(G39) );
  XNOR2_X1 U832 ( .A(G131), .B(n786), .ZN(G33) );
endmodule

