

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717;

  INV_X1 U358 ( .A(G953), .ZN(n710) );
  OR2_X1 U359 ( .A1(n368), .A2(n583), .ZN(n367) );
  NAND2_X2 U360 ( .A1(n372), .A2(n370), .ZN(n584) );
  AND2_X1 U361 ( .A1(n520), .A2(n376), .ZN(n400) );
  XNOR2_X2 U362 ( .A(n401), .B(KEYINPUT32), .ZN(n715) );
  NOR2_X1 U363 ( .A1(n593), .A2(n691), .ZN(n595) );
  NAND2_X1 U364 ( .A1(n558), .A2(n524), .ZN(n634) );
  XNOR2_X2 U365 ( .A(n365), .B(G134), .ZN(n349) );
  XNOR2_X2 U366 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X2 U367 ( .A(G113), .B(G116), .ZN(n395) );
  XNOR2_X1 U368 ( .A(n387), .B(KEYINPUT39), .ZN(n348) );
  NOR2_X1 U369 ( .A1(n529), .A2(n536), .ZN(n505) );
  INV_X1 U370 ( .A(KEYINPUT78), .ZN(n382) );
  NOR2_X1 U371 ( .A1(n583), .A2(n582), .ZN(n618) );
  NAND2_X1 U372 ( .A1(n348), .A2(n571), .ZN(n573) );
  NAND2_X1 U373 ( .A1(n412), .A2(n408), .ZN(n407) );
  AND2_X1 U374 ( .A1(n414), .A2(n413), .ZN(n412) );
  AND2_X1 U375 ( .A1(n374), .A2(n373), .ZN(n372) );
  XNOR2_X1 U376 ( .A(n642), .B(n427), .ZN(n559) );
  NAND2_X2 U377 ( .A1(n362), .A2(n359), .ZN(n642) );
  XNOR2_X1 U378 ( .A(n349), .B(n429), .ZN(n705) );
  XNOR2_X1 U379 ( .A(n514), .B(n338), .ZN(n464) );
  XNOR2_X1 U380 ( .A(n438), .B(n437), .ZN(n704) );
  NAND2_X1 U381 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X1 U382 ( .A(KEYINPUT35), .B(n382), .ZN(n366) );
  NOR2_X2 U383 ( .A1(n521), .A2(n402), .ZN(n401) );
  XNOR2_X2 U384 ( .A(n347), .B(n548), .ZN(n696) );
  NOR2_X1 U385 ( .A1(n634), .A2(n579), .ZN(n540) );
  XNOR2_X2 U386 ( .A(n519), .B(G469), .ZN(n579) );
  XOR2_X1 U387 ( .A(KEYINPUT72), .B(KEYINPUT5), .Z(n450) );
  XOR2_X1 U388 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n438) );
  XNOR2_X1 U389 ( .A(G902), .B(KEYINPUT15), .ZN(n589) );
  AND2_X1 U390 ( .A1(n622), .A2(n388), .ZN(n563) );
  AND2_X1 U391 ( .A1(n577), .A2(n389), .ZN(n388) );
  INV_X1 U392 ( .A(n559), .ZN(n389) );
  OR2_X1 U393 ( .A1(n599), .A2(n360), .ZN(n359) );
  AND2_X1 U394 ( .A1(n364), .A2(n363), .ZN(n362) );
  NAND2_X1 U395 ( .A1(n456), .A2(n361), .ZN(n360) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n486) );
  XOR2_X1 U397 ( .A(KEYINPUT68), .B(G131), .Z(n480) );
  AND2_X1 U398 ( .A1(n355), .A2(n383), .ZN(n354) );
  XNOR2_X1 U399 ( .A(G116), .B(G107), .ZN(n500) );
  INV_X1 U400 ( .A(G143), .ZN(n432) );
  OR2_X1 U401 ( .A1(n635), .A2(n634), .ZN(n537) );
  INV_X1 U402 ( .A(KEYINPUT73), .ZN(n410) );
  XNOR2_X1 U403 ( .A(n579), .B(KEYINPUT1), .ZN(n635) );
  XNOR2_X1 U404 ( .A(n424), .B(n423), .ZN(n422) );
  XNOR2_X1 U405 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U406 ( .A(G119), .B(G110), .ZN(n423) );
  XNOR2_X1 U407 ( .A(n705), .B(n448), .ZN(n517) );
  INV_X1 U408 ( .A(KEYINPUT36), .ZN(n381) );
  XNOR2_X1 U409 ( .A(n527), .B(n528), .ZN(n368) );
  AND2_X1 U410 ( .A1(n665), .A2(n541), .ZN(n527) );
  NAND2_X1 U411 ( .A1(n371), .A2(n337), .ZN(n370) );
  NAND2_X1 U412 ( .A1(n651), .A2(KEYINPUT19), .ZN(n373) );
  XNOR2_X1 U413 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n510) );
  BUF_X1 U414 ( .A(n635), .Z(n386) );
  XNOR2_X1 U415 ( .A(n446), .B(n339), .ZN(n425) );
  OR2_X1 U416 ( .A1(n689), .A2(G902), .ZN(n426) );
  INV_X1 U417 ( .A(KEYINPUT6), .ZN(n427) );
  XNOR2_X1 U418 ( .A(n602), .B(KEYINPUT59), .ZN(n434) );
  OR2_X1 U419 ( .A1(n670), .A2(n343), .ZN(n358) );
  INV_X1 U420 ( .A(G210), .ZN(n369) );
  INV_X1 U421 ( .A(KEYINPUT46), .ZN(n352) );
  NOR2_X1 U422 ( .A1(n654), .A2(n620), .ZN(n586) );
  INV_X1 U423 ( .A(KEYINPUT70), .ZN(n451) );
  XOR2_X1 U424 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n485) );
  XNOR2_X1 U425 ( .A(G104), .B(G122), .ZN(n484) );
  XNOR2_X1 U426 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U427 ( .A(G113), .ZN(n481) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n488) );
  XNOR2_X1 U429 ( .A(KEYINPUT66), .B(G101), .ZN(n470) );
  XNOR2_X1 U430 ( .A(n480), .B(n430), .ZN(n429) );
  XNOR2_X1 U431 ( .A(n431), .B(G137), .ZN(n430) );
  INV_X1 U432 ( .A(KEYINPUT4), .ZN(n431) );
  XOR2_X1 U433 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n467) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n457) );
  XOR2_X1 U435 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n458) );
  OR2_X1 U436 ( .A1(G237), .A2(G902), .ZN(n477) );
  NOR2_X1 U437 ( .A1(n650), .A2(n651), .ZN(n656) );
  INV_X1 U438 ( .A(G902), .ZN(n361) );
  NAND2_X1 U439 ( .A1(n428), .A2(G902), .ZN(n363) );
  NOR2_X1 U440 ( .A1(n633), .A2(n420), .ZN(n419) );
  INV_X1 U441 ( .A(n632), .ZN(n420) );
  INV_X1 U442 ( .A(KEYINPUT45), .ZN(n548) );
  NOR2_X1 U443 ( .A1(n714), .A2(n545), .ZN(n546) );
  XNOR2_X1 U444 ( .A(n393), .B(n391), .ZN(n590) );
  XNOR2_X1 U445 ( .A(n499), .B(n392), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n500), .B(G122), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n512), .B(n511), .ZN(n513) );
  INV_X1 U448 ( .A(KEYINPUT74), .ZN(n511) );
  XNOR2_X1 U449 ( .A(n526), .B(n525), .ZN(n665) );
  INV_X1 U450 ( .A(KEYINPUT33), .ZN(n525) );
  NAND2_X1 U451 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U452 ( .A(n496), .B(n495), .ZN(n535) );
  XNOR2_X1 U453 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U454 ( .A1(G902), .A2(n601), .ZN(n496) );
  INV_X1 U455 ( .A(G475), .ZN(n493) );
  NOR2_X1 U456 ( .A1(n378), .A2(n579), .ZN(n585) );
  XNOR2_X1 U457 ( .A(n578), .B(n379), .ZN(n378) );
  INV_X1 U458 ( .A(KEYINPUT28), .ZN(n379) );
  INV_X1 U459 ( .A(KEYINPUT0), .ZN(n403) );
  NOR2_X1 U460 ( .A1(n536), .A2(n535), .ZN(n571) );
  NAND2_X1 U461 ( .A1(n687), .A2(G472), .ZN(n418) );
  XNOR2_X1 U462 ( .A(n444), .B(n704), .ZN(n689) );
  XNOR2_X1 U463 ( .A(n440), .B(n422), .ZN(n443) );
  XNOR2_X1 U464 ( .A(n590), .B(KEYINPUT124), .ZN(n591) );
  XNOR2_X1 U465 ( .A(n565), .B(n380), .ZN(n566) );
  XNOR2_X1 U466 ( .A(n381), .B(KEYINPUT109), .ZN(n380) );
  OR2_X1 U467 ( .A1(n386), .A2(n558), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n571), .B(n390), .ZN(n622) );
  INV_X1 U469 ( .A(KEYINPUT105), .ZN(n390) );
  NOR2_X1 U470 ( .A1(n433), .A2(n691), .ZN(n605) );
  AND2_X1 U471 ( .A1(n357), .A2(n356), .ZN(n679) );
  XNOR2_X1 U472 ( .A(n358), .B(n678), .ZN(n357) );
  NOR2_X1 U473 ( .A1(n651), .A2(KEYINPUT19), .ZN(n337) );
  XNOR2_X1 U474 ( .A(KEYINPUT16), .B(G122), .ZN(n338) );
  XOR2_X1 U475 ( .A(KEYINPUT88), .B(KEYINPUT25), .Z(n339) );
  AND2_X1 U476 ( .A1(n407), .A2(n415), .ZN(n340) );
  INV_X1 U477 ( .A(n456), .ZN(n428) );
  AND2_X1 U478 ( .A1(n520), .A2(n386), .ZN(n341) );
  XNOR2_X1 U479 ( .A(n642), .B(KEYINPUT104), .ZN(n567) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n558) );
  XOR2_X1 U481 ( .A(n599), .B(n598), .Z(n342) );
  OR2_X1 U482 ( .A1(n589), .A2(n369), .ZN(n343) );
  XNOR2_X1 U483 ( .A(KEYINPUT79), .B(KEYINPUT48), .ZN(n344) );
  XOR2_X1 U484 ( .A(n600), .B(KEYINPUT63), .Z(n345) );
  NOR2_X1 U485 ( .A1(G952), .A2(n710), .ZN(n691) );
  INV_X1 U486 ( .A(n691), .ZN(n356) );
  NAND2_X1 U487 ( .A1(n547), .A2(n546), .ZN(n347) );
  XNOR2_X1 U488 ( .A(n353), .B(n352), .ZN(n351) );
  XNOR2_X1 U489 ( .A(n350), .B(n344), .ZN(n421) );
  NOR2_X4 U490 ( .A1(n670), .A2(n589), .ZN(n687) );
  XNOR2_X2 U491 ( .A(n346), .B(KEYINPUT2), .ZN(n670) );
  NOR2_X2 U492 ( .A1(n696), .A2(n708), .ZN(n346) );
  NAND2_X1 U493 ( .A1(n520), .A2(n559), .ZN(n521) );
  XNOR2_X2 U494 ( .A(n385), .B(n510), .ZN(n520) );
  NAND2_X1 U495 ( .A1(n354), .A2(n351), .ZN(n350) );
  XNOR2_X2 U496 ( .A(n692), .B(n365), .ZN(n377) );
  NAND2_X1 U497 ( .A1(n348), .A2(n588), .ZN(n632) );
  XNOR2_X1 U498 ( .A(n349), .B(n502), .ZN(n393) );
  NAND2_X1 U499 ( .A1(n717), .A2(n405), .ZN(n353) );
  AND2_X1 U500 ( .A1(n436), .A2(n587), .ZN(n355) );
  NAND2_X1 U501 ( .A1(n599), .A2(n428), .ZN(n364) );
  NOR2_X1 U502 ( .A1(n567), .A2(n651), .ZN(n568) );
  XNOR2_X2 U503 ( .A(n447), .B(n432), .ZN(n365) );
  XNOR2_X2 U504 ( .A(n367), .B(n366), .ZN(n716) );
  NAND2_X1 U505 ( .A1(n687), .A2(G478), .ZN(n592) );
  NOR2_X1 U506 ( .A1(n549), .A2(n651), .ZN(n375) );
  INV_X1 U507 ( .A(n549), .ZN(n371) );
  NAND2_X1 U508 ( .A1(n549), .A2(KEYINPUT19), .ZN(n374) );
  NAND2_X1 U509 ( .A1(n564), .A2(n375), .ZN(n565) );
  AND2_X1 U510 ( .A1(n567), .A2(n386), .ZN(n376) );
  XNOR2_X2 U511 ( .A(n377), .B(n474), .ZN(n675) );
  OR2_X1 U512 ( .A1(n716), .A2(KEYINPUT44), .ZN(n531) );
  AND2_X1 U513 ( .A1(n574), .A2(n415), .ZN(n406) );
  NAND2_X1 U514 ( .A1(n687), .A2(G475), .ZN(n435) );
  XNOR2_X1 U515 ( .A(n384), .B(n523), .ZN(n530) );
  XNOR2_X1 U516 ( .A(n435), .B(n434), .ZN(n433) );
  AND2_X2 U517 ( .A1(n399), .A2(n638), .ZN(n613) );
  NOR2_X2 U518 ( .A1(n613), .A2(n715), .ZN(n384) );
  XNOR2_X1 U519 ( .A(n568), .B(KEYINPUT30), .ZN(n415) );
  NAND2_X1 U520 ( .A1(n406), .A2(n407), .ZN(n387) );
  INV_X1 U521 ( .A(n629), .ZN(n383) );
  NAND2_X1 U522 ( .A1(n509), .A2(n541), .ZN(n385) );
  XNOR2_X1 U523 ( .A(n400), .B(KEYINPUT64), .ZN(n399) );
  NAND2_X1 U524 ( .A1(n584), .A2(n479), .ZN(n404) );
  NOR2_X1 U525 ( .A1(n683), .A2(G902), .ZN(n519) );
  XNOR2_X2 U526 ( .A(n394), .B(n453), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n451), .A2(KEYINPUT83), .ZN(n397) );
  NAND2_X1 U528 ( .A1(n452), .A2(KEYINPUT70), .ZN(n398) );
  XNOR2_X2 U529 ( .A(n404), .B(n403), .ZN(n541) );
  XNOR2_X2 U530 ( .A(n465), .B(n464), .ZN(n692) );
  XNOR2_X1 U531 ( .A(n405), .B(G131), .ZN(G33) );
  XNOR2_X2 U532 ( .A(n573), .B(n572), .ZN(n405) );
  OR2_X1 U533 ( .A1(n569), .A2(n409), .ZN(n408) );
  INV_X1 U534 ( .A(n570), .ZN(n411) );
  NAND2_X1 U535 ( .A1(n570), .A2(KEYINPUT73), .ZN(n413) );
  NAND2_X1 U536 ( .A1(n569), .A2(KEYINPUT73), .ZN(n414) );
  XNOR2_X1 U537 ( .A(n416), .B(n345), .ZN(G57) );
  NAND2_X1 U538 ( .A1(n417), .A2(n356), .ZN(n416) );
  XNOR2_X1 U539 ( .A(n418), .B(n342), .ZN(n417) );
  NAND2_X1 U540 ( .A1(n421), .A2(n419), .ZN(n708) );
  NOR2_X2 U541 ( .A1(n537), .A2(n559), .ZN(n526) );
  XNOR2_X2 U542 ( .A(n463), .B(G107), .ZN(n514) );
  XNOR2_X2 U543 ( .A(G110), .B(G104), .ZN(n463) );
  XNOR2_X1 U544 ( .A(n517), .B(n518), .ZN(n683) );
  XNOR2_X1 U545 ( .A(n517), .B(n455), .ZN(n599) );
  XNOR2_X1 U546 ( .A(n618), .B(KEYINPUT77), .ZN(n436) );
  XNOR2_X1 U547 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U548 ( .A(n465), .B(n454), .ZN(n455) );
  XNOR2_X1 U549 ( .A(n704), .B(n483), .ZN(n492) );
  INV_X1 U550 ( .A(KEYINPUT112), .ZN(n600) );
  INV_X1 U551 ( .A(KEYINPUT125), .ZN(n594) );
  XOR2_X1 U552 ( .A(G146), .B(G125), .Z(n469) );
  XNOR2_X1 U553 ( .A(G140), .B(n469), .ZN(n437) );
  XNOR2_X1 U554 ( .A(G137), .B(G128), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n439), .B(KEYINPUT87), .ZN(n440) );
  NAND2_X1 U556 ( .A1(G234), .A2(n710), .ZN(n441) );
  XOR2_X1 U557 ( .A(KEYINPUT8), .B(n441), .Z(n501) );
  NAND2_X1 U558 ( .A1(G221), .A2(n501), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U560 ( .A1(G234), .A2(n589), .ZN(n445) );
  XNOR2_X1 U561 ( .A(KEYINPUT20), .B(n445), .ZN(n506) );
  NAND2_X1 U562 ( .A1(n506), .A2(G217), .ZN(n446) );
  XNOR2_X1 U563 ( .A(G472), .B(KEYINPUT92), .ZN(n456) );
  XNOR2_X2 U564 ( .A(G128), .B(KEYINPUT75), .ZN(n447) );
  XOR2_X1 U565 ( .A(G146), .B(n470), .Z(n448) );
  NAND2_X1 U566 ( .A1(n486), .A2(G210), .ZN(n449) );
  XOR2_X1 U567 ( .A(n450), .B(n449), .Z(n454) );
  INV_X1 U568 ( .A(KEYINPUT83), .ZN(n452) );
  XOR2_X1 U569 ( .A(G119), .B(KEYINPUT3), .Z(n453) );
  INV_X1 U570 ( .A(n567), .ZN(n576) );
  NOR2_X1 U571 ( .A1(G898), .A2(n710), .ZN(n694) );
  XNOR2_X1 U572 ( .A(n458), .B(n457), .ZN(n460) );
  NAND2_X1 U573 ( .A1(n460), .A2(G902), .ZN(n459) );
  XNOR2_X1 U574 ( .A(n459), .B(KEYINPUT85), .ZN(n550) );
  NAND2_X1 U575 ( .A1(n694), .A2(n550), .ZN(n462) );
  NAND2_X1 U576 ( .A1(G952), .A2(n460), .ZN(n664) );
  NOR2_X1 U577 ( .A1(G953), .A2(n664), .ZN(n554) );
  INV_X1 U578 ( .A(n554), .ZN(n461) );
  NAND2_X1 U579 ( .A1(n462), .A2(n461), .ZN(n479) );
  NAND2_X1 U580 ( .A1(G224), .A2(n710), .ZN(n466) );
  XNOR2_X1 U581 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U582 ( .A(n469), .B(n468), .Z(n473) );
  INV_X1 U583 ( .A(n470), .ZN(n471) );
  XNOR2_X1 U584 ( .A(KEYINPUT4), .B(n471), .ZN(n472) );
  XNOR2_X1 U585 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U586 ( .A1(n675), .A2(n589), .ZN(n476) );
  NAND2_X1 U587 ( .A1(G210), .A2(n477), .ZN(n475) );
  XNOR2_X2 U588 ( .A(n476), .B(n475), .ZN(n549) );
  NAND2_X1 U589 ( .A1(G214), .A2(n477), .ZN(n478) );
  XOR2_X1 U590 ( .A(KEYINPUT84), .B(n478), .Z(n651) );
  XNOR2_X1 U591 ( .A(G143), .B(n480), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n490) );
  NAND2_X1 U593 ( .A1(G214), .A2(n486), .ZN(n487) );
  XNOR2_X1 U594 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U595 ( .A(n490), .B(n489), .Z(n491) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n601) );
  XNOR2_X1 U597 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n494) );
  INV_X1 U598 ( .A(n535), .ZN(n529) );
  XNOR2_X1 U599 ( .A(KEYINPUT99), .B(G478), .ZN(n504) );
  XOR2_X1 U600 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n498) );
  XNOR2_X1 U601 ( .A(KEYINPUT98), .B(KEYINPUT9), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U603 ( .A1(G217), .A2(n501), .ZN(n502) );
  NOR2_X1 U604 ( .A1(G902), .A2(n590), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n504), .B(n503), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n505), .B(KEYINPUT102), .ZN(n652) );
  XOR2_X1 U607 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n508) );
  NAND2_X1 U608 ( .A1(n506), .A2(G221), .ZN(n507) );
  XNOR2_X1 U609 ( .A(n508), .B(n507), .ZN(n639) );
  XOR2_X1 U610 ( .A(n639), .B(KEYINPUT90), .Z(n524) );
  AND2_X1 U611 ( .A1(n652), .A2(n524), .ZN(n509) );
  NAND2_X1 U612 ( .A1(G227), .A2(n710), .ZN(n512) );
  XOR2_X1 U613 ( .A(n515), .B(KEYINPUT86), .Z(n516) );
  XNOR2_X1 U614 ( .A(n516), .B(G140), .ZN(n518) );
  INV_X1 U615 ( .A(n558), .ZN(n638) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U617 ( .A1(n522), .A2(KEYINPUT80), .ZN(n523) );
  INV_X1 U618 ( .A(KEYINPUT34), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n536), .A2(n529), .ZN(n583) );
  NAND2_X1 U620 ( .A1(n530), .A2(n716), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n532), .A2(n531), .ZN(n547) );
  AND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n533) );
  NAND2_X1 U623 ( .A1(n341), .A2(n533), .ZN(n534) );
  XNOR2_X1 U624 ( .A(KEYINPUT103), .B(n534), .ZN(n714) );
  NAND2_X1 U625 ( .A1(n536), .A2(n535), .ZN(n615) );
  XOR2_X1 U626 ( .A(KEYINPUT100), .B(n615), .Z(n588) );
  NOR2_X1 U627 ( .A1(n571), .A2(n588), .ZN(n654) );
  XOR2_X1 U628 ( .A(KEYINPUT31), .B(KEYINPUT93), .Z(n539) );
  NOR2_X1 U629 ( .A1(n642), .A2(n537), .ZN(n646) );
  NAND2_X1 U630 ( .A1(n646), .A2(n541), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n627) );
  XNOR2_X1 U632 ( .A(n540), .B(KEYINPUT91), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n642), .A2(n541), .ZN(n542) );
  NOR2_X1 U634 ( .A1(n569), .A2(n542), .ZN(n608) );
  NOR2_X1 U635 ( .A1(n627), .A2(n608), .ZN(n543) );
  NOR2_X1 U636 ( .A1(n654), .A2(n543), .ZN(n544) );
  XOR2_X1 U637 ( .A(KEYINPUT101), .B(n544), .Z(n545) );
  INV_X1 U638 ( .A(n549), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G953), .A2(n550), .ZN(n551) );
  NOR2_X1 U640 ( .A1(G900), .A2(n551), .ZN(n552) );
  XNOR2_X1 U641 ( .A(n552), .B(KEYINPUT106), .ZN(n553) );
  NOR2_X1 U642 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U643 ( .A(KEYINPUT76), .B(n555), .ZN(n570) );
  NOR2_X1 U644 ( .A1(n639), .A2(n570), .ZN(n556) );
  XNOR2_X1 U645 ( .A(n556), .B(KEYINPUT69), .ZN(n557) );
  NOR2_X1 U646 ( .A1(n558), .A2(n557), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n386), .A2(n563), .ZN(n560) );
  NOR2_X1 U648 ( .A1(n651), .A2(n560), .ZN(n561) );
  XNOR2_X1 U649 ( .A(n561), .B(KEYINPUT43), .ZN(n562) );
  NOR2_X1 U650 ( .A1(n581), .A2(n562), .ZN(n633) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(n563), .ZN(n564) );
  NOR2_X1 U652 ( .A1(n386), .A2(n566), .ZN(n629) );
  XOR2_X1 U653 ( .A(KEYINPUT38), .B(n581), .Z(n574) );
  XOR2_X1 U654 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n572) );
  INV_X1 U655 ( .A(n574), .ZN(n650) );
  NAND2_X1 U656 ( .A1(n652), .A2(n656), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n575), .B(KEYINPUT41), .ZN(n666) );
  AND2_X1 U658 ( .A1(n576), .A2(n577), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n666), .A2(n585), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n580), .B(KEYINPUT42), .ZN(n717) );
  NAND2_X1 U661 ( .A1(n581), .A2(n340), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n620) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT47), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n595), .B(n594), .ZN(G63) );
  XOR2_X1 U666 ( .A(KEYINPUT111), .B(KEYINPUT82), .Z(n597) );
  XNOR2_X1 U667 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n597), .B(n596), .ZN(n598) );
  INV_X1 U669 ( .A(n601), .ZN(n602) );
  INV_X1 U670 ( .A(KEYINPUT123), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT60), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n605), .B(n604), .ZN(G60) );
  XOR2_X1 U673 ( .A(G104), .B(KEYINPUT113), .Z(n607) );
  NAND2_X1 U674 ( .A1(n608), .A2(n622), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n607), .B(n606), .ZN(G6) );
  XNOR2_X1 U676 ( .A(G107), .B(KEYINPUT27), .ZN(n612) );
  XOR2_X1 U677 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n610) );
  INV_X1 U678 ( .A(n615), .ZN(n626) );
  NAND2_X1 U679 ( .A1(n608), .A2(n626), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n612), .B(n611), .ZN(G9) );
  BUF_X1 U682 ( .A(n613), .Z(n614) );
  XOR2_X1 U683 ( .A(G110), .B(n614), .Z(G12) );
  NOR2_X1 U684 ( .A1(n615), .A2(n620), .ZN(n617) );
  XNOR2_X1 U685 ( .A(G128), .B(KEYINPUT29), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n617), .B(n616), .ZN(G30) );
  XOR2_X1 U687 ( .A(G143), .B(n618), .Z(G45) );
  INV_X1 U688 ( .A(n622), .ZN(n619) );
  NOR2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U690 ( .A(G146), .B(n621), .Z(G48) );
  XOR2_X1 U691 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n624) );
  NAND2_X1 U692 ( .A1(n627), .A2(n622), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U694 ( .A(G113), .B(n625), .ZN(G15) );
  NAND2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(G116), .ZN(G18) );
  XNOR2_X1 U697 ( .A(G125), .B(n629), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U699 ( .A(G134), .B(KEYINPUT117), .Z(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(G36) );
  XOR2_X1 U701 ( .A(G140), .B(n633), .Z(G42) );
  XOR2_X1 U702 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n637) );
  NAND2_X1 U703 ( .A1(n386), .A2(n634), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(n644) );
  NAND2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U706 ( .A(KEYINPUT49), .B(n640), .Z(n641) );
  NAND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U710 ( .A(n647), .B(KEYINPUT119), .Z(n648) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(n648), .ZN(n649) );
  NAND2_X1 U712 ( .A1(n666), .A2(n649), .ZN(n661) );
  NAND2_X1 U713 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U714 ( .A1(n653), .A2(n652), .ZN(n658) );
  INV_X1 U715 ( .A(n654), .ZN(n655) );
  NAND2_X1 U716 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U717 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U718 ( .A1(n665), .A2(n659), .ZN(n660) );
  NAND2_X1 U719 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U720 ( .A(KEYINPUT52), .B(n662), .Z(n663) );
  NOR2_X1 U721 ( .A1(n664), .A2(n663), .ZN(n669) );
  NAND2_X1 U722 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U723 ( .A(KEYINPUT120), .B(n667), .Z(n668) );
  NOR2_X1 U724 ( .A1(n669), .A2(n668), .ZN(n672) );
  BUF_X1 U725 ( .A(n670), .Z(n671) );
  NAND2_X1 U726 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U727 ( .A1(n673), .A2(G953), .ZN(n674) );
  XNOR2_X1 U728 ( .A(n674), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U729 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n677) );
  XNOR2_X1 U730 ( .A(n675), .B(KEYINPUT81), .ZN(n676) );
  XNOR2_X1 U731 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U732 ( .A(KEYINPUT56), .B(n679), .ZN(G51) );
  XOR2_X1 U733 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n681) );
  XNOR2_X1 U734 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n680) );
  XNOR2_X1 U735 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U736 ( .A(n683), .B(n682), .Z(n685) );
  NAND2_X1 U737 ( .A1(n687), .A2(G469), .ZN(n684) );
  XNOR2_X1 U738 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n691), .A2(n686), .ZN(G54) );
  NAND2_X1 U740 ( .A1(G217), .A2(n687), .ZN(n688) );
  XNOR2_X1 U741 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U742 ( .A1(n691), .A2(n690), .ZN(G66) );
  XOR2_X1 U743 ( .A(n692), .B(G101), .Z(n693) );
  NOR2_X1 U744 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U745 ( .A(KEYINPUT127), .B(n695), .Z(n703) );
  NOR2_X1 U746 ( .A1(G953), .A2(n696), .ZN(n697) );
  XOR2_X1 U747 ( .A(KEYINPUT126), .B(n697), .Z(n701) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n698) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n698), .ZN(n699) );
  NAND2_X1 U750 ( .A1(n699), .A2(G898), .ZN(n700) );
  NAND2_X1 U751 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(G69) );
  XNOR2_X1 U753 ( .A(n705), .B(n704), .ZN(n709) );
  XNOR2_X1 U754 ( .A(G227), .B(n709), .ZN(n706) );
  NAND2_X1 U755 ( .A1(G900), .A2(n706), .ZN(n707) );
  NAND2_X1 U756 ( .A1(n707), .A2(G953), .ZN(n713) );
  XNOR2_X1 U757 ( .A(n709), .B(n708), .ZN(n711) );
  NAND2_X1 U758 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U759 ( .A1(n713), .A2(n712), .ZN(G72) );
  XOR2_X1 U760 ( .A(G101), .B(n714), .Z(G3) );
  XOR2_X1 U761 ( .A(n715), .B(G119), .Z(G21) );
  XNOR2_X1 U762 ( .A(G122), .B(n716), .ZN(G24) );
  XNOR2_X1 U763 ( .A(G137), .B(n717), .ZN(G39) );
endmodule

