//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(G234), .A2(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G952), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT21), .B(G898), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(G902), .A3(G953), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G210), .B1(G237), .B2(G902), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT5), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G116), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(G113), .B(new_n201), .C1(new_n203), .C2(new_n199), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT2), .B(G113), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n213), .A2(KEYINPUT78), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(G104), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n225));
  AOI211_X1 g039(.A(new_n225), .B(new_n222), .C1(new_n216), .C2(new_n219), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n207), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(G110), .B(G122), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n216), .B2(new_n219), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n209), .A2(new_n212), .A3(new_n215), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(new_n205), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n206), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n227), .A2(new_n229), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n227), .A2(KEYINPUT84), .A3(new_n239), .A4(new_n229), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT6), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n227), .A2(new_n239), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n228), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n229), .B(new_n247), .C1(new_n227), .C2(new_n239), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n252), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n260), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(G146), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n262), .A2(new_n267), .A3(G125), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT1), .B1(new_n266), .B2(new_n256), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(G128), .B1(new_n258), .B2(new_n257), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n264), .B(new_n273), .C1(new_n266), .C2(new_n256), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n269), .B1(G125), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n189), .A2(G224), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT85), .Z(new_n279));
  XNOR2_X1  g093(.A(new_n277), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n251), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n217), .A2(new_n218), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n217), .A2(new_n218), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n223), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n207), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n207), .A2(new_n285), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n228), .B(KEYINPUT8), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n276), .A2(G125), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT7), .B(new_n278), .C1(new_n290), .C2(new_n268), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n269), .B(new_n292), .C1(G125), .C2(new_n276), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n289), .B(new_n294), .C1(new_n242), .C2(new_n243), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n198), .B1(new_n282), .B2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n245), .A2(new_n228), .B1(KEYINPUT83), .B2(KEYINPUT6), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(new_n249), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n280), .B1(new_n299), .B2(new_n244), .ZN(new_n300));
  INV_X1    g114(.A(new_n198), .ZN(new_n301));
  NOR4_X1   g115(.A1(new_n300), .A2(new_n295), .A3(G902), .A4(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n187), .B(new_n197), .C1(new_n297), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  AND4_X1   g119(.A1(G143), .A2(new_n305), .A3(new_n189), .A4(G214), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  AOI21_X1  g121(.A(G143), .B1(new_n307), .B2(G214), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n189), .A3(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n256), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT87), .A3(G131), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(KEYINPUT17), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT89), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT75), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n252), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n320), .A2(G146), .A3(new_n323), .A4(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n306), .A2(new_n308), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT87), .B1(new_n315), .B2(G131), .ZN(new_n338));
  AOI211_X1 g152(.A(new_n310), .B(new_n336), .C1(new_n313), .C2(new_n314), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n334), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n311), .A2(new_n316), .A3(new_n341), .A4(KEYINPUT17), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n318), .A2(new_n333), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n253), .A2(new_n255), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n319), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n321), .A2(G125), .ZN(new_n346));
  OAI21_X1  g160(.A(G146), .B1(new_n325), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n313), .A2(new_n314), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT18), .B(G131), .C1(new_n306), .C2(new_n308), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT86), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n335), .A2(new_n349), .B1(new_n345), .B2(new_n347), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n352), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n343), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n208), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT90), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n304), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n343), .A2(new_n358), .A3(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(G475), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n343), .A2(new_n361), .A3(new_n358), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT19), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n319), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT19), .B1(new_n325), .B2(new_n346), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n344), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n331), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n367), .B(new_n361), .C1(new_n358), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n356), .B1(new_n355), .B2(new_n352), .ZN(new_n377));
  AND4_X1   g191(.A1(new_n356), .A2(new_n352), .A3(new_n348), .A4(new_n350), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n315), .A2(G131), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n311), .B2(new_n316), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n377), .A2(new_n378), .B1(new_n380), .B2(new_n373), .ZN(new_n381));
  INV_X1    g195(.A(new_n361), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT88), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n366), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n365), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G116), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(G116), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT93), .ZN(new_n396));
  INV_X1    g210(.A(new_n393), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  OAI21_X1  g212(.A(G107), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n397), .A2(new_n392), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n211), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n256), .B2(G128), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n272), .A2(KEYINPUT92), .A3(G143), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n403), .A2(new_n404), .B1(G128), .B2(new_n256), .ZN(new_n405));
  INV_X1    g219(.A(G134), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n400), .B(new_n211), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n404), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(G134), .A3(new_n405), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n405), .B1(new_n412), .B2(G134), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT9), .B(G234), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT71), .B(G217), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n418), .A2(G953), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT94), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n415), .A3(new_n421), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(KEYINPUT94), .A3(new_n422), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n304), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n428), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(new_n365), .C1(new_n387), .C2(new_n388), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n390), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n263), .B1(new_n344), .B2(G143), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n272), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n274), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n220), .A2(new_n223), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n270), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n259), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n274), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n222), .B1(new_n216), .B2(new_n219), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G137), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G134), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT11), .B1(new_n406), .B2(G137), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n445), .A3(G134), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n446), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(KEYINPUT65), .A3(new_n336), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n336), .A2(KEYINPUT65), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n452), .B(new_n446), .C1(new_n447), .C2(new_n449), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n444), .A2(KEYINPUT12), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n285), .A2(new_n225), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n441), .B2(new_n274), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n262), .A2(new_n267), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n237), .B1(new_n231), .B2(new_n233), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n463), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n469));
  AOI211_X1 g283(.A(KEYINPUT80), .B(new_n469), .C1(new_n443), .C2(new_n438), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n471));
  INV_X1    g285(.A(new_n469), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n439), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n454), .B(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n468), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n189), .A2(G227), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  AND3_X1   g293(.A1(new_n460), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n439), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT80), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n465), .B1(new_n224), .B2(new_n226), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n466), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n439), .A2(new_n471), .A3(new_n472), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n455), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n479), .B1(new_n487), .B2(new_n476), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n435), .B(new_n304), .C1(new_n480), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n475), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n444), .A2(KEYINPUT12), .A3(new_n455), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n444), .B2(new_n455), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n486), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n479), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n476), .A3(new_n479), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(G469), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(G469), .A2(G902), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G221), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n417), .B2(new_n304), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n303), .A2(new_n434), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT24), .B(G110), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n272), .A2(G119), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n200), .A2(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n272), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT73), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(KEYINPUT23), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n516), .A3(KEYINPUT23), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n508), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n511), .B1(new_n519), .B2(G110), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n331), .A3(new_n345), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(G110), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n332), .C1(new_n510), .C2(new_n507), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n526), .B(KEYINPUT76), .Z(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n521), .B2(new_n523), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n304), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT25), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n420), .B1(G234), .B2(new_n304), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT25), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n304), .C1(new_n527), .C2(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n532), .A4(new_n534), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n527), .A2(new_n529), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n532), .A2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n543));
  OR3_X1    g357(.A1(new_n445), .A2(KEYINPUT66), .A3(G134), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n445), .A2(G134), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT66), .B1(new_n445), .B2(G134), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n544), .A2(G131), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n450), .B2(G131), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n271), .B2(new_n275), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n262), .B(new_n267), .C1(new_n451), .C2(new_n453), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n236), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n236), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT68), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n307), .A2(G210), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n558), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n549), .A2(new_n551), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n236), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n568), .B2(new_n556), .ZN(new_n569));
  INV_X1    g383(.A(new_n556), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT28), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n554), .A2(new_n573), .A3(new_n556), .A4(new_n563), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G472), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n304), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT69), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .A4(new_n304), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(KEYINPUT69), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n569), .A2(new_n571), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT29), .B1(new_n585), .B2(new_n563), .ZN(new_n586));
  INV_X1    g400(.A(new_n554), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n562), .B1(new_n587), .B2(new_n570), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(KEYINPUT29), .A3(new_n563), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n543), .B1(new_n584), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n576), .B1(new_n589), .B2(new_n590), .ZN(new_n594));
  AOI211_X1 g408(.A(KEYINPUT70), .B(new_n594), .C1(new_n582), .C2(new_n583), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n504), .B(new_n542), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  AND3_X1   g411(.A1(new_n575), .A2(new_n576), .A3(new_n304), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n576), .B1(new_n575), .B2(new_n304), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n542), .A2(new_n600), .A3(new_n502), .A4(new_n499), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT95), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n390), .A2(new_n433), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n426), .A2(new_n604), .A3(new_n427), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n416), .B2(new_n422), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT96), .B(new_n421), .C1(new_n408), .C2(new_n415), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT33), .B(new_n425), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n605), .A2(new_n609), .A3(G478), .A4(new_n304), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n428), .A2(new_n429), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n602), .A2(new_n303), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n618), .A2(KEYINPUT97), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n357), .A2(new_n354), .B1(new_n368), .B2(new_n374), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n367), .B1(new_n620), .B2(new_n361), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n381), .A2(KEYINPUT88), .A3(new_n382), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n359), .A2(new_n361), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n386), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT20), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n618), .A2(KEYINPUT97), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n619), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n428), .B(new_n430), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n365), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n617), .B1(new_n303), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n187), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n251), .A2(new_n281), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n304), .A3(new_n296), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n301), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n282), .A2(new_n198), .A3(new_n296), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n629), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(KEYINPUT98), .A3(new_n637), .A4(new_n197), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n602), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G107), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  AND2_X1   g456(.A1(new_n521), .A2(new_n523), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n645), .B2(new_n647), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n540), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n537), .A3(new_n538), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n187), .B(new_n651), .C1(new_n297), .C2(new_n302), .ZN(new_n652));
  INV_X1    g466(.A(new_n599), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n499), .A2(new_n577), .A3(new_n653), .A4(new_n502), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n652), .A2(new_n654), .A3(new_n434), .A4(new_n196), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n584), .A2(new_n592), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT70), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n584), .A2(new_n543), .A3(new_n592), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n503), .ZN(new_n662));
  INV_X1    g476(.A(new_n652), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n191), .B1(new_n195), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n629), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n662), .A3(new_n663), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  AOI21_X1  g482(.A(new_n563), .B1(new_n568), .B2(new_n556), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n587), .A2(new_n570), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n670), .B2(new_n563), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n584), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n651), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n634), .A2(new_n635), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n634), .A2(KEYINPUT38), .A3(new_n635), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n665), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n662), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n499), .A2(new_n684), .A3(new_n502), .A4(new_n681), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n431), .B1(new_n390), .B2(new_n433), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n187), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n675), .A2(new_n680), .A3(new_n683), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  INV_X1    g503(.A(new_n665), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n625), .A2(new_n618), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n432), .B1(new_n691), .B2(new_n365), .ZN(new_n692));
  INV_X1    g506(.A(new_n433), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n612), .B(new_n690), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n603), .A2(new_n696), .A3(new_n612), .A4(new_n690), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n661), .A2(new_n662), .A3(new_n699), .A4(new_n663), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NOR2_X1   g515(.A1(new_n303), .A2(new_n613), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n480), .A2(new_n488), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n304), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n502), .A3(new_n489), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n661), .A2(new_n542), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND2_X1  g524(.A1(new_n638), .A2(new_n630), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n661), .A2(new_n711), .A3(new_n542), .A4(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NOR3_X1   g527(.A1(new_n652), .A2(new_n434), .A3(new_n196), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n661), .A2(new_n714), .A3(new_n707), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n686), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n676), .A2(new_n187), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n603), .B2(new_n628), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n600), .A2(KEYINPUT102), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(KEYINPUT102), .B2(new_n653), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(new_n542), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n197), .A3(new_n724), .A4(new_n707), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n651), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n719), .A2(new_n706), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n699), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NAND3_X1  g545(.A1(new_n634), .A2(new_n187), .A3(new_n635), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n695), .A2(new_n697), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n592), .A2(new_n579), .A3(new_n581), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n542), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(KEYINPUT104), .A3(new_n662), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n695), .A2(new_n733), .A3(new_n662), .A4(new_n697), .ZN(new_n741));
  INV_X1    g555(.A(new_n736), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n732), .A2(new_n503), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n542), .B(new_n746), .C1(new_n593), .C2(new_n595), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n737), .B1(new_n747), .B2(new_n698), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n748), .A3(KEYINPUT105), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n661), .A2(new_n542), .A3(new_n666), .A4(new_n746), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n650), .A2(new_n537), .A3(new_n538), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n600), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n390), .A2(new_n761), .A3(new_n433), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n761), .B1(new_n390), .B2(new_n433), .ZN(new_n763));
  OAI211_X1 g577(.A(KEYINPUT43), .B(new_n612), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n390), .B(new_n433), .C1(KEYINPUT108), .C2(new_n612), .ZN(new_n766));
  INV_X1    g580(.A(new_n612), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n757), .B(new_n760), .C1(new_n764), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT110), .B1(new_n771), .B2(new_n732), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT106), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n495), .B2(new_n496), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(new_n435), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n479), .B1(new_n486), .B2(new_n490), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n454), .B1(new_n468), .B2(new_n474), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n479), .B1(new_n460), .B2(new_n476), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT106), .A3(G469), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n496), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n775), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n498), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT107), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n498), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n489), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n791), .A3(new_n786), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(new_n502), .A3(new_n681), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n764), .A2(new_n770), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n759), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n757), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(KEYINPUT44), .A3(new_n759), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n733), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n772), .A2(new_n794), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  AOI21_X1  g616(.A(KEYINPUT47), .B1(new_n793), .B2(new_n502), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n793), .A2(KEYINPUT47), .A3(new_n502), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n593), .A2(new_n595), .ZN(new_n807));
  INV_X1    g621(.A(new_n542), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n734), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(G952), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n189), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n767), .B1(new_n692), .B2(new_n693), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n434), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n601), .A3(new_n303), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n655), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n596), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n596), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n732), .A2(new_n758), .A3(new_n665), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n627), .A2(new_n431), .A3(new_n365), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n661), .A2(new_n662), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n662), .A2(new_n695), .A3(new_n697), .A4(new_n733), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT113), .B1(new_n828), .B2(new_n728), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n741), .A2(new_n830), .A3(new_n727), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n755), .B(new_n827), .C1(new_n829), .C2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n708), .A2(new_n712), .A3(new_n715), .A4(new_n725), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n824), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n758), .A2(new_n502), .A3(new_n499), .A4(new_n690), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT114), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n721), .A3(new_n673), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n667), .A2(new_n700), .A3(new_n730), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n503), .B1(new_n659), .B2(new_n660), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n663), .C1(new_n666), .C2(new_n699), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n730), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n834), .A2(new_n753), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n834), .A2(new_n844), .A3(KEYINPUT53), .A4(new_n749), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n834), .A2(new_n753), .A3(new_n844), .A4(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n847), .A2(new_n855), .A3(new_n848), .A4(new_n849), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n705), .A2(new_n501), .A3(new_n489), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n804), .A2(new_n805), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n190), .B1(new_n764), .B2(new_n770), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n724), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n733), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n862), .B2(KEYINPUT117), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n706), .A2(new_n732), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n674), .A2(new_n542), .A3(new_n191), .A4(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n603), .A3(new_n612), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n187), .B(new_n706), .C1(new_n678), .C2(new_n679), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n860), .A3(new_n724), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT50), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n866), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n860), .A2(new_n864), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n728), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n862), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n863), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT48), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n876), .A2(new_n742), .B1(KEYINPUT118), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(KEYINPUT118), .B2(new_n880), .ZN(new_n882));
  OR4_X1    g696(.A1(KEYINPUT118), .A2(new_n875), .A3(new_n880), .A4(new_n736), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n814), .B(G953), .C1(new_n861), .C2(new_n729), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n863), .B2(new_n878), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n865), .A2(new_n613), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n879), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n815), .B1(new_n857), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n705), .A2(new_n489), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n542), .B1(new_n890), .B2(KEYINPUT49), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(KEYINPUT49), .B2(new_n890), .ZN(new_n892));
  INV_X1    g706(.A(new_n680), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n612), .B1(new_n762), .B2(new_n763), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n501), .A3(new_n631), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .A4(new_n674), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n889), .A2(new_n896), .ZN(G75));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n304), .C1(new_n847), .C2(new_n849), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n251), .A2(new_n281), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n300), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n899), .A2(KEYINPUT56), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n304), .B1(new_n847), .B2(new_n849), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G210), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n189), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(G51));
  XOR2_X1   g724(.A(new_n498), .B(KEYINPUT57), .Z(new_n911));
  AND3_X1   g725(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n703), .ZN(new_n915));
  INV_X1    g729(.A(new_n784), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n905), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n909), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n909), .B1(new_n919), .B2(new_n623), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .A4(new_n384), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT58), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n923), .B(new_n304), .C1(new_n847), .C2(new_n849), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(G475), .A4(new_n384), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n920), .A2(new_n922), .A3(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(new_n605), .A2(new_n609), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n912), .B2(new_n913), .ZN(new_n932));
  INV_X1    g746(.A(new_n909), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n930), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n857), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n936), .B2(new_n928), .ZN(G63));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n938), .B(new_n939), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n847), .B2(new_n849), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(new_n539), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n648), .B2(new_n649), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n933), .A4(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n933), .B1(new_n942), .B2(new_n539), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n648), .A2(new_n649), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n948), .B(new_n941), .C1(new_n847), .C2(new_n849), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n950), .ZN(G66));
  INV_X1    g765(.A(G224), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n193), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n824), .A2(new_n833), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(G953), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n299), .B(new_n244), .C1(G898), .C2(new_n189), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n667), .A2(new_n700), .A3(new_n688), .A4(new_n730), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n842), .A2(KEYINPUT62), .A3(new_n688), .A4(new_n730), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n961), .A2(new_n962), .B1(new_n806), .B2(new_n811), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n807), .A2(new_n808), .A3(new_n682), .A4(new_n817), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n733), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n801), .A2(KEYINPUT122), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT122), .B1(new_n801), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n189), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n552), .A2(new_n553), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT121), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n370), .A2(new_n371), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n958), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  AOI211_X1 g789(.A(KEYINPUT123), .B(new_n973), .C1(new_n968), .C2(new_n189), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n794), .A2(new_n721), .A3(new_n742), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n753), .A2(new_n812), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n842), .A2(new_n730), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n801), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n801), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n980), .A2(new_n986), .A3(new_n189), .A4(new_n755), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n973), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n977), .B(new_n989), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n772), .A2(new_n800), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n797), .A2(new_n502), .A3(new_n681), .A4(new_n793), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n965), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT122), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n801), .A2(KEYINPUT122), .A3(new_n965), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n1000), .B2(new_n963), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT123), .B1(new_n1001), .B2(new_n973), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n969), .A2(new_n958), .A3(new_n974), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n989), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n990), .A3(new_n1003), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n991), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n993), .A2(new_n1006), .ZN(G72));
  XNOR2_X1  g821(.A(new_n670), .B(KEYINPUT126), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n755), .A2(new_n980), .A3(new_n986), .A4(new_n954), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n562), .B(new_n1008), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n847), .B2(new_n852), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n588), .A2(new_n564), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n909), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n963), .B(new_n954), .C1(new_n966), .C2(new_n967), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1008), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1018), .A2(KEYINPUT127), .A3(new_n563), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT127), .B1(new_n1018), .B2(new_n563), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1013), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(G57));
endmodule


