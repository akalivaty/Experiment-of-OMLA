//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n195), .C1(G119), .C2(new_n194), .ZN(new_n196));
  XNOR2_X1  g010(.A(G119), .B(G128), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT24), .B(G110), .Z(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n205), .A3(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(KEYINPUT72), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n199), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n196), .A2(G110), .B1(new_n197), .B2(new_n198), .ZN(new_n214));
  XNOR2_X1  g028(.A(G125), .B(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n209), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n190), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G902), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n217), .A3(new_n190), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT74), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(KEYINPUT74), .B2(new_n223), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G234), .B2(new_n220), .ZN(new_n228));
  INV_X1    g042(.A(new_n221), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n229), .A2(new_n218), .A3(G902), .ZN(new_n230));
  INV_X1    g044(.A(new_n224), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n226), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(new_n218), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n228), .A2(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT31), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n238), .B(new_n243), .C1(new_n239), .C2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G134), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n242), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n239), .A2(G137), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n249), .B2(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n207), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  AND4_X1   g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .A4(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n194), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n255), .B2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT66), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n258), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n252), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n261), .B1(new_n259), .B2(new_n260), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(KEYINPUT66), .A3(new_n265), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n257), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n272), .B2(new_n251), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n241), .A2(new_n244), .A3(new_n247), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n248), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT0), .A4(G128), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n260), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT30), .A4(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT2), .A2(G113), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT2), .A2(G113), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT2), .A3(G113), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G116), .B(G119), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n288), .B1(new_n291), .B2(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n248), .A2(KEYINPUT65), .A3(new_n250), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT65), .B1(new_n248), .B2(new_n250), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n267), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT67), .B(new_n267), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n281), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n296), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n276), .B2(new_n280), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n273), .A3(new_n269), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G210), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G101), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n237), .B1(new_n305), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n296), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n303), .A2(new_n281), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n251), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n248), .A2(KEYINPUT65), .A3(new_n250), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT67), .B1(new_n322), .B2(new_n267), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n297), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n315), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(KEYINPUT31), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n252), .A2(new_n267), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n306), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n306), .A2(new_n273), .A3(new_n269), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n304), .B2(new_n295), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n316), .A2(new_n327), .B1(new_n334), .B2(new_n313), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT32), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n295), .B1(new_n318), .B2(new_n323), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n333), .B1(new_n339), .B2(new_n307), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n313), .B1(new_n340), .B2(new_n329), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT31), .B1(new_n325), .B2(new_n326), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n237), .B(new_n315), .C1(new_n317), .C2(new_n324), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n336), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n269), .A2(new_n273), .A3(new_n281), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n295), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n307), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n329), .B1(new_n350), .B2(KEYINPUT28), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n313), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n334), .A2(new_n313), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n331), .B1(new_n317), .B2(new_n324), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n314), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G472), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n236), .B1(new_n347), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(G104), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT76), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n364), .A2(KEYINPUT76), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n361), .B2(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(new_n367), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n361), .A3(G104), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n367), .A2(KEYINPUT79), .A3(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n272), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n253), .B1(G143), .B2(new_n207), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n194), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n263), .A2(KEYINPUT80), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n260), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n374), .B(new_n382), .C1(new_n389), .C2(new_n257), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n276), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT12), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n276), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT10), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n373), .B1(new_n366), .B2(new_n372), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n399));
  AOI21_X1  g213(.A(new_n279), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n367), .A2(G107), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n368), .B2(new_n370), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n363), .B1(new_n365), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G101), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n374), .A3(KEYINPUT4), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n397), .A2(new_n267), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n254), .A2(new_n386), .A3(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n388), .A2(G128), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n257), .B1(new_n411), .B2(new_n265), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n408), .B(new_n409), .C1(new_n383), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n408), .B1(new_n390), .B2(new_n409), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n395), .B(new_n407), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n405), .A2(new_n374), .A3(KEYINPUT4), .ZN(new_n419));
  OAI211_X1 g233(.A(G101), .B(new_n399), .C1(new_n402), .C2(new_n404), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n280), .A2(new_n420), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n419), .A2(new_n421), .B1(new_n272), .B2(new_n396), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n383), .A2(new_n412), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT81), .B1(new_n423), .B2(KEYINPUT10), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT82), .B1(new_n425), .B2(new_n395), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n394), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n188), .A2(G227), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n416), .A2(new_n417), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n413), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n395), .A4(new_n407), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n425), .A2(new_n395), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n427), .A2(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G469), .B1(new_n436), .B2(G902), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(G469), .C1(new_n436), .C2(G902), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT84), .B(G469), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n433), .ZN(new_n442));
  INV_X1    g256(.A(new_n430), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n442), .A2(new_n394), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n442), .B2(new_n435), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n220), .B(new_n441), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n438), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT9), .B(G234), .ZN(new_n448));
  OAI21_X1  g262(.A(G221), .B1(new_n448), .B2(G902), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT75), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n255), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT90), .A2(G143), .ZN(new_n455));
  OAI211_X1 g269(.A(G214), .B(new_n309), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n309), .A2(G214), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n453), .B2(new_n255), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n458), .A3(new_n242), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G146), .B1(new_n204), .B2(new_n205), .ZN(new_n464));
  INV_X1    g278(.A(new_n209), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT72), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(KEYINPUT17), .A3(G131), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n463), .A2(new_n211), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G113), .B(G122), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n367), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT18), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n456), .B(new_n458), .C1(new_n472), .C2(new_n242), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n215), .B(new_n207), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n473), .B(new_n474), .C1(new_n460), .C2(new_n472), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n471), .B1(new_n469), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n220), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G475), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n215), .B(KEYINPUT19), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n465), .B1(new_n481), .B2(new_n207), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n460), .A2(new_n462), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n475), .ZN(new_n485));
  INV_X1    g299(.A(new_n471), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n490), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT20), .B(new_n492), .C1(new_n487), .C2(new_n488), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n479), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n448), .A2(new_n227), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G116), .ZN(new_n497));
  INV_X1    g311(.A(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G122), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G107), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n499), .A3(new_n361), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n194), .B2(G143), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n255), .A2(KEYINPUT13), .A3(G128), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n194), .A2(G143), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G134), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n194), .A2(G143), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n255), .A2(G128), .ZN(new_n511));
  OR3_X1    g325(.A1(new_n510), .A2(new_n511), .A3(G134), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n514));
  INV_X1    g328(.A(new_n502), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n515), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n498), .A2(KEYINPUT14), .A3(G122), .ZN(new_n518));
  OAI211_X1 g332(.A(G107), .B(new_n518), .C1(new_n500), .C2(KEYINPUT14), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n513), .A2(new_n514), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n503), .A2(KEYINPUT91), .A3(new_n512), .A4(new_n509), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n495), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n495), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT92), .B(new_n220), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n524), .A3(new_n521), .ZN(new_n530));
  INV_X1    g344(.A(new_n495), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n521), .A3(new_n495), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n528), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(KEYINPUT92), .A3(new_n220), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n188), .A2(G952), .ZN(new_n538));
  INV_X1    g352(.A(G234), .ZN(new_n539));
  INV_X1    g353(.A(G237), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n220), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT21), .B(G898), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n494), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n288), .A2(new_n290), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n192), .A2(G116), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n549), .B(G113), .C1(KEYINPUT5), .C2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(KEYINPUT88), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n547), .A2(KEYINPUT88), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n548), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n383), .B2(KEYINPUT88), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n552), .B(new_n554), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n406), .A2(new_n295), .A3(new_n420), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(new_n374), .A3(new_n382), .A4(new_n548), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n553), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n272), .A2(new_n202), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n279), .A2(G125), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT86), .B(G224), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G953), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n558), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n566), .ZN(new_n570));
  INV_X1    g384(.A(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n562), .A2(new_n571), .A3(new_n563), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n567), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  OAI21_X1  g390(.A(G210), .B1(G237), .B2(G902), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n559), .A2(new_n560), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n553), .A2(KEYINPUT85), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n561), .A2(KEYINPUT6), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(KEYINPUT6), .A3(new_n580), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n577), .A3(new_n584), .ZN(new_n586));
  INV_X1    g400(.A(new_n577), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n561), .A2(KEYINPUT6), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n580), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n590), .A2(new_n582), .B1(new_n570), .B2(new_n572), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n558), .A2(new_n561), .A3(new_n568), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n220), .B1(new_n592), .B2(new_n573), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n587), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n594), .A3(KEYINPUT89), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n452), .A2(new_n546), .A3(new_n585), .A4(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n360), .A2(new_n447), .A3(new_n451), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  AND2_X1   g412(.A1(new_n447), .A2(new_n451), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n344), .B2(new_n220), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n335), .A2(new_n337), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(new_n602), .A3(new_n236), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n527), .A2(G902), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n534), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT33), .B1(new_n534), .B2(KEYINPUT93), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n534), .A2(new_n220), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n527), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n545), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n494), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n452), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n586), .B2(new_n594), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(KEYINPUT94), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n586), .A2(new_n594), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n452), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n599), .A2(new_n603), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n491), .A2(new_n493), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n478), .A2(new_n627), .A3(G475), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n478), .B2(G475), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n626), .B(new_n537), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n625), .B1(new_n631), .B2(new_n545), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n491), .A2(new_n493), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n479), .A2(KEYINPUT95), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n628), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(KEYINPUT96), .A3(new_n611), .A4(new_n537), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n599), .A2(new_n603), .A3(new_n615), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT97), .Z(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT35), .B(G107), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NAND2_X1  g455(.A1(new_n213), .A2(new_n217), .ZN(new_n642));
  INV_X1    g456(.A(new_n190), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n234), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n232), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n601), .A2(new_n602), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n447), .A2(new_n451), .A3(new_n596), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NAND2_X1  g466(.A1(new_n615), .A2(new_n647), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n542), .B1(new_n543), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n653), .A2(new_n631), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n335), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n345), .B1(new_n344), .B2(new_n336), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n359), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n447), .A2(new_n656), .A3(new_n659), .A4(new_n451), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n655), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n599), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n599), .A2(new_n666), .A3(new_n662), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n595), .A2(new_n585), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT38), .Z(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n356), .A2(new_n313), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n220), .B1(new_n350), .B2(new_n314), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n347), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n614), .B1(new_n529), .B2(new_n536), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n494), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n647), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT98), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n671), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n665), .B1(new_n664), .B2(new_n667), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  INV_X1    g499(.A(new_n655), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n610), .A2(new_n494), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n653), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n447), .A2(new_n659), .A3(new_n451), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  OAI21_X1  g504(.A(new_n435), .B1(new_n418), .B2(new_n426), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n691), .A2(new_n430), .B1(new_n434), .B2(new_n394), .ZN(new_n692));
  OAI21_X1  g506(.A(G469), .B1(new_n692), .B2(G902), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n449), .A3(new_n446), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n360), .A2(new_n621), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT41), .B(G113), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT100), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n696), .B(new_n698), .ZN(G15));
  AND4_X1   g513(.A1(new_n449), .A2(new_n693), .A3(new_n446), .A4(new_n615), .ZN(new_n700));
  INV_X1    g514(.A(new_n236), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n659), .A3(new_n701), .A4(new_n637), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  INV_X1    g517(.A(new_n653), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n695), .A2(new_n659), .A3(new_n546), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  AND2_X1   g520(.A1(new_n586), .A2(new_n594), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT101), .B1(new_n707), .B2(new_n678), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n618), .A2(new_n709), .A3(new_n494), .A4(new_n677), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n545), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n316), .A2(new_n327), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n351), .A2(new_n314), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n337), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n601), .A2(new_n236), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n695), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NOR4_X1   g531(.A1(new_n601), .A2(new_n714), .A3(new_n687), .A4(new_n648), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n700), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  INV_X1    g535(.A(new_n449), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n437), .B2(new_n446), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n614), .B1(new_n595), .B2(new_n585), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n659), .A2(new_n723), .A3(new_n701), .A4(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n721), .B1(new_n725), .B2(new_n687), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n427), .A2(new_n430), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n434), .A2(new_n435), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(G469), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n446), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n731), .A2(new_n449), .A3(new_n724), .ZN(new_n732));
  INV_X1    g546(.A(new_n687), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n360), .A3(KEYINPUT42), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NOR2_X1   g550(.A1(new_n631), .A2(new_n655), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n360), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n647), .B1(new_n601), .B2(new_n602), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT104), .Z(new_n742));
  AND2_X1   g556(.A1(new_n607), .A2(new_n609), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(KEYINPUT43), .A3(new_n494), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n494), .A2(new_n745), .B1(new_n609), .B2(new_n607), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n745), .B2(new_n494), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n747), .B2(KEYINPUT43), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n740), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n724), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n727), .A2(new_n728), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n436), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n446), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT102), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n759), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n449), .B(new_n662), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n742), .A2(new_n740), .A3(new_n749), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n751), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n245), .ZN(G39));
  INV_X1    g582(.A(new_n724), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n659), .A2(new_n769), .A3(new_n701), .A4(new_n687), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n449), .B1(new_n762), .B2(new_n764), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(KEYINPUT47), .B(new_n449), .C1(new_n762), .C2(new_n764), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n200), .ZN(G42));
  AND4_X1   g591(.A1(new_n696), .A2(new_n702), .A3(new_n705), .A4(new_n716), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n634), .A2(new_n628), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n537), .A2(new_n655), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n626), .A2(new_n779), .A3(new_n647), .A4(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n724), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n447), .A2(new_n782), .A3(new_n659), .A4(new_n451), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n732), .A2(new_n718), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n738), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n778), .A2(new_n785), .A3(new_n735), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n669), .A2(new_n612), .A3(new_n614), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n447), .A2(new_n451), .A3(new_n603), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n597), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n787), .B1(new_n597), .B2(new_n789), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n447), .A2(new_n451), .A3(new_n603), .ZN(new_n792));
  INV_X1    g606(.A(new_n537), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n494), .A2(new_n793), .A3(new_n545), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n452), .A3(new_n595), .A4(new_n585), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT107), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n650), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n790), .A2(new_n791), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n786), .A2(new_n798), .A3(KEYINPUT108), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n597), .A2(new_n789), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT106), .ZN(new_n802));
  INV_X1    g616(.A(new_n797), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n597), .A2(new_n787), .A3(new_n789), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n778), .A2(new_n785), .A3(new_n735), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n648), .A2(new_n686), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n708), .B2(new_n710), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n675), .A3(new_n723), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT109), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n675), .A3(new_n813), .A4(new_n723), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n660), .A2(new_n689), .A3(new_n719), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n808), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n660), .A2(new_n689), .A3(new_n719), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n812), .A2(new_n814), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n799), .A2(new_n807), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n798), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n778), .A2(KEYINPUT112), .A3(new_n735), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n778), .B2(new_n735), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n817), .A2(new_n832), .A3(new_n820), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n828), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n825), .A4(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n799), .A2(new_n807), .A3(new_n821), .ZN(new_n837));
  INV_X1    g651(.A(new_n823), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n799), .A2(new_n807), .A3(new_n834), .A4(new_n833), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n837), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n841), .B2(new_n825), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n834), .A2(new_n833), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n827), .A2(new_n830), .A3(new_n829), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n843), .A2(new_n844), .B1(new_n822), .B2(new_n823), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT113), .B1(new_n845), .B2(new_n825), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n824), .A2(new_n835), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n839), .A2(new_n840), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n799), .A2(new_n807), .A3(new_n821), .A4(new_n838), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n854), .A3(new_n855), .A4(new_n836), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n694), .A2(new_n769), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n748), .A2(new_n542), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n748), .A2(new_n862), .A3(new_n542), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT48), .A4(new_n360), .ZN(new_n865));
  INV_X1    g679(.A(new_n715), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n861), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n700), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n675), .A2(new_n236), .A3(new_n541), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n858), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n610), .A2(new_n494), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n872), .A3(new_n538), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(new_n360), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n865), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n610), .A2(new_n494), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n601), .A2(new_n648), .A3(new_n714), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n879), .B2(new_n864), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n670), .A2(new_n694), .A3(new_n452), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT50), .B1(new_n867), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n693), .A2(new_n450), .A3(new_n446), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n774), .A2(new_n775), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n867), .A2(new_n724), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n876), .B1(new_n889), .B2(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n891), .B(new_n884), .C1(new_n886), .C2(new_n888), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT118), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n886), .A2(new_n888), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n889), .A2(KEYINPUT51), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n876), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n847), .A2(new_n856), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT119), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n847), .A2(new_n899), .A3(new_n856), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT120), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  OR4_X1    g720(.A1(new_n236), .A2(new_n747), .A3(new_n450), .A4(new_n614), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT105), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n670), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n693), .A2(new_n446), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT49), .Z(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n910), .A3(new_n676), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(G75));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n581), .A2(new_n583), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n578), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n845), .A2(new_n220), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G210), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n915), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n921), .B2(new_n920), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n188), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n918), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n849), .B(KEYINPUT54), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n757), .B(KEYINPUT57), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n445), .B2(new_n444), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n845), .A2(new_n220), .A3(new_n756), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(G54));
  AND3_X1   g748(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n935), .B2(new_n489), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n935), .B2(new_n489), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n935), .A2(KEYINPUT122), .A3(new_n489), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(G60));
  OR2_X1    g754(.A1(new_n605), .A2(new_n606), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n847), .A2(new_n856), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n929), .A2(new_n941), .A3(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n924), .A3(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n845), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n925), .B1(new_n950), .B2(new_n233), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n645), .B2(new_n950), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n565), .B2(new_n544), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n798), .A2(new_n778), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n916), .B1(G898), .B2(new_n188), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  AOI21_X1  g773(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n324), .A2(new_n282), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n481), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n188), .A2(G900), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n735), .A2(new_n738), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n708), .A2(new_n710), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n360), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n965), .B(new_n818), .C1(new_n765), .C2(new_n967), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n776), .A2(new_n767), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(G953), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT124), .B(new_n964), .C1(new_n969), .C2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n962), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n684), .A2(new_n977), .A3(new_n818), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n776), .A2(new_n767), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n818), .B1(new_n682), .B2(new_n683), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n626), .A2(new_n479), .A3(new_n537), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n769), .B1(new_n871), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n664), .A2(new_n360), .A3(new_n667), .A4(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n978), .A2(new_n979), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n985), .B2(new_n188), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT126), .B(new_n960), .C1(new_n975), .C2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n972), .B2(new_n973), .ZN(new_n989));
  INV_X1    g803(.A(new_n960), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n986), .A2(KEYINPUT123), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT123), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n994), .B(new_n976), .C1(new_n985), .C2(new_n188), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n974), .B(new_n990), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n969), .B2(new_n956), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n356), .A2(new_n313), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n925), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n356), .B2(new_n314), .ZN(new_n1008));
  OAI211_X1 g822(.A(KEYINPUT127), .B(new_n313), .C1(new_n305), .C2(new_n331), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1008), .B(new_n1009), .C1(new_n305), .C2(new_n315), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n853), .A2(new_n1002), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1002), .B1(new_n985), .B2(new_n955), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1006), .B(new_n1011), .C1(new_n672), .C2(new_n1012), .ZN(G57));
endmodule


