//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n203), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n206), .B(new_n217), .C1(new_n220), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G50), .B(G68), .Z(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n218), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n219), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G150), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n219), .A2(new_n247), .ZN(new_n248));
  OAI22_X1  g0048(.A1(new_n244), .A2(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n219), .B1(new_n221), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n243), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n243), .B1(new_n253), .B2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n252), .B(new_n255), .C1(G50), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT9), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n259), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G222), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n265), .B1(new_n266), .B2(new_n263), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n247), .C2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n272), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n277), .B2(G226), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT67), .B(G200), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n271), .A2(G190), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT10), .B1(new_n262), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n261), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n260), .B(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT10), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(new_n282), .A4(new_n281), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(new_n257), .C1(G179), .C2(new_n279), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n274), .B1(new_n277), .B2(G244), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT65), .Z(new_n294));
  INV_X1    g0094(.A(G107), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n267), .A2(new_n211), .B1(new_n295), .B2(new_n263), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n300), .A2(new_n209), .A3(G1698), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n270), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n280), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n244), .A2(new_n248), .B1(new_n219), .B2(new_n266), .ZN(new_n305));
  OR2_X1    g0105(.A1(KEYINPUT15), .A2(G87), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT15), .A2(G87), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n245), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n243), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(new_n310), .B(KEYINPUT66), .Z(new_n311));
  NOR2_X1   g0111(.A1(new_n256), .A2(G77), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n254), .B2(G77), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n304), .B(new_n315), .C1(new_n316), .C2(new_n303), .ZN(new_n317));
  INV_X1    g0117(.A(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n303), .A2(new_n290), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(G179), .C2(new_n303), .ZN(new_n320));
  AND4_X1   g0120(.A1(new_n289), .A2(new_n292), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n276), .A2(new_n272), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n322), .A2(new_n211), .B1(new_n273), .B2(new_n272), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n267), .B2(new_n209), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n263), .A2(KEYINPUT69), .A3(G232), .A4(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n323), .B1(new_n329), .B2(new_n270), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI211_X1 g0132(.A(KEYINPUT13), .B(new_n323), .C1(new_n329), .C2(new_n270), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(G179), .B1(new_n335), .B2(KEYINPUT14), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n334), .A2(new_n290), .B1(new_n335), .B2(KEYINPUT14), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(KEYINPUT14), .ZN(new_n338));
  OAI211_X1 g0138(.A(G169), .B(new_n338), .C1(new_n332), .C2(new_n333), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n256), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n210), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  INV_X1    g0143(.A(new_n254), .ZN(new_n344));
  INV_X1    g0144(.A(new_n243), .ZN(new_n345));
  INV_X1    g0145(.A(new_n245), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G20), .A2(G33), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n348), .A2(KEYINPUT70), .B1(G50), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n353));
  OAI221_X1 g0153(.A(new_n343), .B1(new_n210), .B2(new_n344), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n340), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n334), .A2(G190), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n356), .C1(new_n360), .C2(new_n334), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT74), .ZN(new_n362));
  INV_X1    g0162(.A(G159), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n248), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n350), .A2(KEYINPUT74), .A3(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n208), .A2(new_n210), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n367), .B2(new_n221), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n300), .A2(new_n219), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT7), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G68), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT7), .A2(G20), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n263), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n369), .B(KEYINPUT16), .C1(new_n372), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT75), .B1(new_n247), .B2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n298), .A3(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n297), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n263), .B2(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n210), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n366), .A2(new_n368), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n380), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n379), .A2(new_n391), .A3(new_n243), .ZN(new_n392));
  INV_X1    g0192(.A(new_n244), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n344), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n244), .A2(new_n256), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n263), .A2(G226), .A3(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n263), .A2(G223), .A3(new_n264), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n270), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n274), .B1(new_n277), .B2(G232), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G169), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(G179), .A3(new_n403), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n316), .A2(KEYINPUT76), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n316), .A2(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n402), .A2(new_n415), .A3(new_n403), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n360), .B1(new_n402), .B2(new_n403), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n392), .A3(new_n396), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n263), .A2(new_n376), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n373), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n210), .B1(new_n370), .B2(KEYINPUT7), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n390), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n345), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n418), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n410), .A2(new_n411), .B1(new_n420), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n321), .A2(new_n358), .A3(new_n361), .A4(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n297), .A2(new_n299), .A3(G244), .A4(new_n264), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT4), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(KEYINPUT77), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n297), .A2(new_n299), .A3(G250), .A4(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G283), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n270), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G41), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(G274), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n276), .ZN(new_n449));
  INV_X1    g0249(.A(G257), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n441), .A2(G179), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n440), .B2(new_n270), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n290), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n295), .B1(new_n387), .B2(new_n388), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n350), .A2(G77), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n295), .A2(KEYINPUT6), .A3(G97), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT6), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n239), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n460), .B2(new_n219), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n243), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n256), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n253), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n256), .A2(new_n464), .A3(new_n218), .A4(new_n242), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(G97), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n454), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n468), .B1(new_n473), .B2(G200), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n454), .A2(G190), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n455), .A2(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT86), .B1(new_n478), .B2(KEYINPUT85), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n300), .A2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(G87), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT86), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(KEYINPUT22), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n263), .A2(new_n483), .A3(new_n219), .A4(new_n479), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n219), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n295), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n477), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n479), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n263), .A2(new_n219), .ZN(new_n495));
  INV_X1    g0295(.A(new_n483), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT24), .A3(new_n485), .A4(new_n491), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n243), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n341), .A2(KEYINPUT25), .A3(new_n295), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT25), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n256), .B2(G107), .ZN(new_n502));
  AOI22_X1  g0302(.A1(G107), .A2(new_n466), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n448), .A2(G264), .A3(new_n276), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n448), .A2(KEYINPUT87), .A3(G264), .A4(new_n276), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n263), .A2(G250), .A3(new_n264), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n263), .A2(G257), .A3(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n506), .A2(new_n507), .B1(new_n511), .B2(new_n270), .ZN(new_n512));
  AOI21_X1  g0312(.A(G200), .B1(new_n512), .B2(new_n447), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n511), .A2(new_n270), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n504), .A2(new_n447), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n514), .A2(G190), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n499), .B(new_n503), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n253), .A2(G45), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n518), .A2(G250), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n276), .B1(G274), .B2(new_n443), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n297), .A2(new_n299), .A3(G244), .A4(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n297), .A2(new_n299), .A3(G238), .A4(new_n264), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n486), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n276), .B1(new_n524), .B2(KEYINPUT79), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n522), .A2(new_n523), .A3(new_n526), .A4(new_n486), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n521), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n280), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n466), .A2(G87), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n219), .B1(new_n326), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G97), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n481), .A2(new_n535), .A3(new_n295), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n297), .A2(new_n299), .A3(new_n219), .A4(G68), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n533), .B1(new_n245), .B2(new_n535), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n243), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n256), .B1(new_n306), .B2(new_n307), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n532), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(KEYINPUT80), .B(new_n542), .C1(new_n540), .C2(new_n243), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n531), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n530), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n528), .A2(G190), .ZN(new_n548));
  AOI211_X1 g0348(.A(G179), .B(new_n521), .C1(new_n525), .C2(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n524), .A2(KEYINPUT79), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n270), .A3(new_n527), .ZN(new_n551));
  AOI21_X1  g0351(.A(G169), .B1(new_n551), .B2(new_n520), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n308), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n466), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n544), .B2(new_n545), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n547), .A2(new_n548), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n476), .A2(new_n517), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n297), .A2(new_n299), .A3(G257), .A4(new_n264), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n297), .A2(new_n299), .A3(G264), .A4(G1698), .ZN(new_n560));
  INV_X1    g0360(.A(G303), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n263), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n270), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n448), .A2(G270), .A3(new_n276), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(new_n447), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n563), .A2(new_n565), .A3(G179), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n256), .A2(new_n464), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT81), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n345), .A4(G116), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT81), .B1(new_n465), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n438), .B(new_n219), .C1(G33), .C2(new_n535), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(G20), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n243), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n243), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n253), .A2(new_n571), .A3(G13), .A4(G20), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT82), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n566), .A2(new_n567), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n567), .B1(new_n566), .B2(new_n583), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n563), .A2(new_n565), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT21), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n290), .B1(KEYINPUT83), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n583), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(KEYINPUT83), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n583), .A2(new_n587), .A3(new_n591), .A4(new_n589), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n514), .B2(new_n515), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n506), .A2(new_n507), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n511), .A2(new_n270), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(G179), .A4(new_n447), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n499), .A2(new_n503), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n586), .B(new_n595), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n583), .B1(G200), .B2(new_n587), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n563), .A2(new_n565), .A3(new_n415), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NOR4_X1   g0409(.A1(new_n431), .A2(new_n558), .A3(new_n605), .A4(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n420), .A2(new_n429), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n361), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n358), .B2(new_n320), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n410), .A2(new_n411), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n289), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n292), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n462), .A2(new_n467), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n475), .B(new_n619), .C1(new_n360), .C2(new_n454), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n462), .A2(new_n470), .A3(new_n467), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n470), .B1(new_n462), .B2(new_n467), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n290), .B1(new_n441), .B2(new_n452), .ZN(new_n624));
  INV_X1    g0424(.A(G179), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n625), .B(new_n451), .C1(new_n440), .C2(new_n270), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n620), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n551), .A2(new_n520), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n280), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n542), .B1(new_n540), .B2(new_n243), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(new_n532), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n632), .A3(new_n548), .A4(new_n531), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n290), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n528), .A2(new_n625), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n556), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n517), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n593), .B(new_n594), .C1(new_n584), .C2(new_n585), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT89), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT89), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n600), .A2(new_n601), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n638), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n636), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n633), .A2(new_n472), .A3(new_n455), .A4(new_n636), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n468), .B1(new_n624), .B2(new_n626), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT90), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n455), .A2(new_n653), .A3(new_n468), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n557), .A2(new_n651), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n648), .B2(new_n655), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n645), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n618), .B1(new_n431), .B2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n253), .A2(new_n219), .A3(G13), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(KEYINPUT92), .A3(KEYINPUT27), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT92), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n664));
  OAI221_X1 g0464(.A(G213), .B1(KEYINPUT27), .B2(new_n661), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n583), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n609), .B1(new_n639), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n642), .B2(new_n668), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n603), .A2(new_n604), .ZN(new_n673));
  INV_X1    g0473(.A(new_n517), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n601), .A2(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n667), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n643), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n667), .B1(new_n586), .B2(new_n595), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n675), .A2(new_n681), .B1(new_n644), .B2(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n204), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n536), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n224), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT96), .ZN(new_n691));
  INV_X1    g0491(.A(new_n604), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n639), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n691), .B1(new_n558), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n638), .A2(new_n605), .A3(KEYINPUT96), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n557), .A2(new_n654), .A3(new_n651), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n646), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n678), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n658), .A2(new_n704), .A3(new_n678), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n638), .A2(new_n694), .A3(new_n608), .A4(new_n678), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT95), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n673), .A2(new_n639), .A3(new_n609), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT95), .A3(new_n638), .A4(new_n678), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n566), .A2(KEYINPUT93), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n587), .B2(new_n625), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n454), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n528), .A2(new_n512), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n512), .A2(new_n447), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(new_n625), .A3(new_n587), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(KEYINPUT94), .A3(new_n473), .A4(new_n629), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n715), .A2(new_n454), .ZN(new_n722));
  INV_X1    g0522(.A(new_n717), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n723), .A4(new_n713), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT94), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n719), .A2(new_n629), .A3(new_n625), .A4(new_n587), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n454), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n718), .A2(new_n721), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n667), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n718), .B(new_n724), .C1(new_n454), .C2(new_n726), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n709), .A2(new_n711), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n706), .B1(G330), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n690), .B1(new_n739), .B2(G1), .ZN(G364));
  OR2_X1    g0540(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n670), .A2(new_n671), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n253), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n685), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n741), .B2(new_n742), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n218), .B1(G20), .B2(new_n290), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n280), .A2(G20), .A3(new_n625), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(new_n316), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n752), .A2(new_n755), .B1(new_n757), .B2(new_n561), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G20), .A3(new_n316), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n263), .B1(new_n761), .B2(G329), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n219), .A2(new_n625), .A3(new_n360), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n316), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n415), .A2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(G326), .ZN(new_n768));
  INV_X1    g0568(.A(G294), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n219), .B1(new_n759), .B2(G190), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n758), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT99), .B1(G20), .B2(G179), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(KEYINPUT99), .A2(G20), .A3(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(new_n316), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n415), .A2(new_n776), .A3(new_n775), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n772), .B1(new_n773), .B2(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT102), .Z(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n300), .B1(new_n785), .B2(G50), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n755), .A2(new_n295), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n760), .A2(new_n363), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n756), .A2(G87), .ZN(new_n791));
  AND4_X1   g0591(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n764), .A2(new_n210), .B1(new_n535), .B2(new_n770), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT101), .Z(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n266), .C2(new_n777), .ZN(new_n795));
  INV_X1    g0595(.A(new_n781), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(G58), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n751), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n748), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n684), .A2(new_n300), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n571), .B2(new_n684), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n421), .A2(new_n422), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n684), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n224), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n237), .A2(new_n442), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n751), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n799), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n670), .B2(new_n809), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n750), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n648), .A2(new_n655), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT91), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n648), .A2(new_n655), .A3(new_n649), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n667), .B1(new_n819), .B2(new_n645), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n318), .A2(new_n667), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n317), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n320), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n320), .A2(new_n667), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n820), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n734), .A2(G330), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n748), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n751), .A2(new_n807), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n799), .B1(new_n266), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n751), .ZN(new_n833));
  INV_X1    g0633(.A(new_n764), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n785), .A2(G137), .B1(new_n834), .B2(G150), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n363), .B2(new_n777), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n796), .B2(G143), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n802), .B1(new_n839), .B2(new_n760), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n754), .A2(G68), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n757), .B2(new_n250), .ZN(new_n842));
  INV_X1    g0642(.A(new_n770), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n840), .B(new_n842), .C1(G58), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n796), .A2(G294), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n300), .B1(new_n760), .B2(new_n773), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n767), .A2(new_n561), .B1(new_n764), .B2(new_n752), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G97), .C2(new_n843), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n754), .A2(G87), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(new_n295), .C2(new_n757), .ZN(new_n851));
  INV_X1    g0651(.A(new_n777), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(G116), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n838), .A2(new_n845), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n832), .B1(new_n833), .B2(new_n854), .C1(new_n826), .C2(new_n808), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n830), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n460), .ZN(new_n857));
  OAI211_X1 g0657(.A(G116), .B(new_n220), .C1(new_n857), .C2(KEYINPUT35), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(KEYINPUT35), .B2(new_n857), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n861));
  OAI21_X1  g0661(.A(G77), .B1(new_n208), .B2(new_n210), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n224), .A2(new_n862), .B1(G50), .B2(new_n210), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n744), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT104), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  INV_X1    g0667(.A(new_n665), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n397), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n419), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT105), .B1(new_n397), .B2(new_n407), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n397), .A2(new_n407), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT37), .B1(new_n873), .B2(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n426), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n425), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n396), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n405), .A2(new_n406), .A3(new_n665), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n419), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n868), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n883), .B(KEYINPUT38), .C1(new_n430), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n874), .A2(new_n872), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n614), .B2(new_n611), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n867), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n430), .B2(new_n869), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n614), .A2(new_n611), .ZN(new_n894));
  INV_X1    g0694(.A(new_n869), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n870), .B2(new_n873), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n875), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n886), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n885), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n891), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n340), .A2(new_n357), .A3(new_n678), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n902), .A2(new_n904), .B1(new_n615), .B2(new_n665), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n357), .A2(new_n667), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n358), .A2(new_n361), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n340), .A2(new_n357), .A3(new_n667), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n658), .A2(new_n678), .A3(new_n826), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n824), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n885), .A2(new_n889), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n709), .A2(new_n711), .A3(new_n731), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n825), .B1(new_n907), .B2(new_n908), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n916), .A3(new_n917), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n921), .A3(G330), .ZN(new_n922));
  INV_X1    g0722(.A(new_n431), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G330), .A3(new_n916), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n918), .A2(new_n921), .A3(new_n923), .A4(new_n916), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n914), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT107), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n704), .B1(new_n701), .B2(new_n678), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n820), .B2(new_n704), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n931), .B2(new_n431), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n923), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n617), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n253), .B2(new_n745), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n928), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n866), .B1(new_n937), .B2(new_n938), .ZN(G367));
  OAI21_X1  g0739(.A(new_n476), .B1(new_n619), .B2(new_n678), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n455), .A2(new_n468), .A3(new_n667), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n682), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT44), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n682), .A2(new_n942), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT45), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n680), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n680), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT111), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(KEYINPUT111), .A3(new_n680), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n675), .A2(new_n681), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n679), .B2(new_n681), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(new_n672), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n738), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n685), .B(KEYINPUT41), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n746), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n672), .A2(new_n679), .A3(new_n942), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n546), .A2(new_n667), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n557), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n636), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT110), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n962), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n954), .A2(new_n940), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  AOI22_X1  g0771(.A1(new_n942), .A2(new_n673), .B1(new_n455), .B2(new_n472), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n667), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n969), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n968), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n961), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n803), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n810), .B1(new_n204), .B2(new_n308), .C1(new_n977), .C2(new_n233), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n748), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n764), .A2(new_n769), .B1(new_n295), .B2(new_n770), .ZN(new_n980));
  INV_X1    g0780(.A(new_n802), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n982), .B2(new_n760), .C1(new_n755), .C2(new_n535), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(G311), .C2(new_n785), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n757), .A2(new_n571), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n985), .A2(KEYINPUT46), .B1(new_n752), .B2(new_n777), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(KEYINPUT46), .B2(new_n985), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n984), .B(new_n987), .C1(new_n561), .C2(new_n781), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n208), .A2(new_n757), .B1(new_n755), .B2(new_n266), .ZN(new_n989));
  INV_X1    g0789(.A(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n263), .B1(new_n990), .B2(new_n760), .C1(new_n764), .C2(new_n363), .ZN(new_n991));
  INV_X1    g0791(.A(G143), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n767), .A2(new_n992), .B1(new_n210), .B2(new_n770), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n250), .B2(new_n777), .C1(new_n246), .C2(new_n781), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT47), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n833), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n988), .A2(new_n995), .A3(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n979), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n809), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n965), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n976), .A2(new_n1001), .ZN(G387));
  NOR2_X1   g0802(.A1(new_n738), .A2(new_n956), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n738), .A2(new_n956), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n685), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n977), .B1(new_n230), .B2(G45), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n687), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n800), .ZN(new_n1009));
  AOI21_X1  g0809(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n393), .A2(new_n250), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n687), .B(new_n1010), .C1(new_n1011), .C2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n204), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n799), .B1(new_n1014), .B2(new_n810), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n679), .B2(new_n1000), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n802), .B1(G326), .B2(new_n761), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n781), .A2(new_n982), .B1(new_n561), .B2(new_n777), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT113), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n773), .B2(new_n764), .C1(new_n782), .C2(new_n767), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT48), .Z(new_n1021));
  OAI22_X1  g0821(.A1(new_n757), .A2(new_n769), .B1(new_n752), .B2(new_n770), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1017), .B1(new_n571), .B2(new_n755), .C1(new_n1023), .C2(KEYINPUT49), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n843), .A2(new_n554), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n781), .B2(new_n250), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT112), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n266), .A2(new_n757), .B1(new_n755), .B2(new_n535), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n802), .B1(new_n246), .B2(new_n760), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n767), .A2(new_n363), .B1(new_n764), .B2(new_n244), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1030), .B(new_n1034), .C1(new_n210), .C2(new_n777), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1024), .A2(new_n1025), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1016), .B1(new_n1036), .B2(new_n751), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n747), .B2(new_n957), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1006), .A2(new_n1038), .ZN(G393));
  AOI21_X1  g0839(.A(new_n686), .B1(new_n1003), .B2(new_n953), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n948), .B(KEYINPUT114), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n951), .A2(new_n952), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1043), .B2(new_n1003), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n747), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n834), .A2(G303), .B1(G116), .B2(new_n843), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n769), .B2(new_n777), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT116), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n756), .A2(G283), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n263), .B1(new_n761), .B2(G322), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n788), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n781), .A2(new_n773), .B1(new_n982), .B2(new_n767), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n781), .A2(new_n363), .B1(new_n246), .B2(new_n767), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  NOR2_X1   g0855(.A1(new_n770), .A2(new_n266), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n834), .B2(G50), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n244), .B2(new_n777), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n981), .B1(G143), .B2(new_n761), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n850), .C1(new_n210), .C2(new_n757), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n1060), .B2(KEYINPUT115), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT115), .B2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1051), .A2(new_n1053), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n833), .B1(new_n1063), .B2(KEYINPUT117), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(KEYINPUT117), .B2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n803), .A2(new_n240), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n751), .B(new_n809), .C1(G97), .C2(new_n684), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n799), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1065), .B(new_n1068), .C1(new_n1000), .C2(new_n942), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1044), .A2(new_n1045), .A3(new_n1069), .ZN(G390));
  NOR3_X1   g0870(.A1(new_n887), .A2(new_n888), .A3(new_n886), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n899), .B2(new_n886), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n890), .B1(new_n1072), .B2(new_n867), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n911), .B2(new_n904), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n701), .A2(new_n678), .A3(new_n823), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(new_n824), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n903), .B(new_n901), .C1(new_n1076), .C2(new_n909), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n917), .A2(new_n734), .A3(G330), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT118), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n917), .A2(new_n916), .A3(new_n1080), .A4(G330), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n917), .A2(new_n916), .A3(G330), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT118), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1074), .A2(new_n1077), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT107), .B1(new_n706), .B2(new_n923), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n929), .B(new_n431), .C1(new_n703), .C2(new_n705), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n618), .B(new_n924), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n734), .A2(G330), .A3(new_n826), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n909), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1083), .A2(new_n1089), .A3(new_n1081), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n824), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n820), .B2(new_n826), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1078), .A2(new_n824), .A3(new_n1075), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n916), .A2(G330), .A3(new_n826), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n909), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1090), .A2(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1079), .A2(new_n1084), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT120), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n686), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n934), .A3(new_n924), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n901), .A2(new_n903), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n909), .B1(new_n1075), .B2(new_n824), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n903), .B1(new_n1092), .B2(new_n909), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n1073), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1083), .A2(new_n1081), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1104), .A2(KEYINPUT120), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT119), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1104), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT119), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1100), .B(new_n1113), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n799), .B1(new_n244), .B2(new_n831), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n777), .A2(new_n535), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n785), .A2(G283), .B1(new_n834), .B2(G107), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n263), .B(new_n1056), .C1(G294), .C2(new_n761), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n791), .A3(new_n1123), .A4(new_n841), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(G116), .C2(new_n796), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n781), .A2(new_n839), .B1(new_n1126), .B2(new_n767), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT121), .Z(new_n1128));
  AOI21_X1  g0928(.A(new_n300), .B1(new_n761), .B2(G125), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n363), .B2(new_n770), .C1(new_n990), .C2(new_n764), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n246), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  NAND2_X1  g0932(.A1(new_n852), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT53), .B1(new_n757), .B2(new_n246), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1130), .B(new_n1135), .C1(G50), .C2(new_n754), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1125), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1120), .B1(new_n1137), .B2(new_n833), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1073), .B2(new_n807), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1116), .B2(new_n747), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1119), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(new_n1087), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n289), .A2(new_n292), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n257), .A2(new_n868), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(KEYINPUT124), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(new_n922), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n922), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n914), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n905), .A2(new_n913), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n1151), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1143), .A2(KEYINPUT57), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1114), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT119), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1087), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1165), .A3(new_n685), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1148), .A2(new_n807), .A3(new_n1149), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n250), .B1(G33), .B2(G41), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n981), .B2(new_n275), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n770), .A2(new_n210), .B1(new_n760), .B2(new_n752), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n767), .A2(new_n571), .B1(new_n764), .B2(new_n535), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n554), .C2(new_n852), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n981), .B(new_n275), .C1(new_n757), .C2(new_n266), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n755), .A2(new_n208), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(new_n295), .C2(new_n781), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n785), .A2(G125), .B1(new_n834), .B2(G132), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n246), .B2(new_n770), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n756), .B2(new_n1132), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n1126), .B2(new_n781), .C1(new_n990), .C2(new_n777), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n754), .A2(G159), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n751), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT122), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(KEYINPUT122), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n831), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n748), .B1(new_n1192), .B2(G50), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT123), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1190), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1158), .A2(new_n747), .B1(new_n1167), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1166), .A2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1104), .A2(new_n959), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n300), .B1(new_n760), .B2(new_n561), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n554), .B2(new_n843), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n757), .B2(new_n535), .C1(new_n266), .C2(new_n755), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n785), .A2(G294), .B1(new_n834), .B2(G116), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n295), .B2(new_n777), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1205), .B2(new_n1204), .C1(new_n752), .C2(new_n781), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n802), .B1(new_n1126), .B2(new_n760), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n1174), .C1(G159), .C2(new_n756), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n834), .A2(new_n1132), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n250), .B2(new_n770), .C1(new_n839), .C2(new_n767), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G150), .B2(new_n852), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1209), .B(new_n1212), .C1(new_n990), .C2(new_n781), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n748), .B1(G68), .B2(new_n1192), .C1(new_n1214), .C2(new_n833), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n909), .B2(new_n807), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1103), .B2(new_n747), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1199), .A2(new_n1217), .ZN(G381));
  OR4_X1    g1018(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1196), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1164), .B1(new_n1221), .B2(new_n1142), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n686), .B1(new_n1222), .B2(KEYINPUT57), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1220), .B1(new_n1223), .B2(new_n1165), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G387), .A2(new_n1219), .A3(G381), .A4(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1226), .ZN(G409));
  NAND4_X1  g1028(.A1(G387), .A2(new_n1044), .A3(new_n1045), .A4(new_n1069), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G390), .A2(new_n1001), .A3(new_n976), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(G393), .B(new_n814), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1198), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n1097), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n685), .A3(new_n1104), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1217), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n830), .A3(new_n855), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(G384), .A3(new_n1217), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n666), .A2(G213), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1119), .A2(new_n1140), .A3(new_n1196), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1222), .A2(new_n959), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1246), .B(new_n1250), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT63), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(G2897), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1245), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT63), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1237), .B(new_n1253), .C1(new_n1258), .C2(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1246), .A4(new_n1250), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1260), .A2(new_n1257), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT127), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1260), .A3(new_n1269), .A4(new_n1263), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1259), .B1(new_n1267), .B2(new_n1272), .ZN(G405));
  NAND2_X1  g1073(.A1(new_n1226), .A2(new_n1261), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1246), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1226), .A2(new_n1261), .A3(new_n1245), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(new_n1271), .Z(G402));
endmodule


