

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731;

  NOR2_X1 U374 ( .A1(n550), .A2(n665), .ZN(n386) );
  OR2_X1 U375 ( .A1(n666), .A2(n582), .ZN(n416) );
  NAND2_X1 U376 ( .A1(n580), .A2(n365), .ZN(n420) );
  NOR2_X1 U377 ( .A1(n546), .A2(n544), .ZN(n522) );
  XNOR2_X1 U378 ( .A(n514), .B(n513), .ZN(n546) );
  XNOR2_X1 U379 ( .A(n351), .B(n713), .ZN(n512) );
  XNOR2_X1 U380 ( .A(n506), .B(n361), .ZN(n351) );
  XNOR2_X1 U381 ( .A(n371), .B(n444), .ZN(n532) );
  XNOR2_X1 U382 ( .A(n352), .B(G146), .ZN(n526) );
  INV_X1 U383 ( .A(G125), .ZN(n352) );
  BUF_X1 U384 ( .A(G116), .Z(n425) );
  NOR2_X1 U385 ( .A1(n716), .A2(n355), .ZN(n601) );
  XNOR2_X2 U386 ( .A(n422), .B(n600), .ZN(n716) );
  AND2_X2 U387 ( .A1(n387), .A2(n639), .ZN(n553) );
  XNOR2_X2 U388 ( .A(n540), .B(n388), .ZN(n387) );
  XNOR2_X2 U389 ( .A(n353), .B(n374), .ZN(n680) );
  XNOR2_X2 U390 ( .A(n699), .B(n534), .ZN(n353) );
  XNOR2_X1 U391 ( .A(n526), .B(n453), .ZN(n713) );
  NOR2_X1 U392 ( .A1(n639), .A2(n638), .ZN(n547) );
  XOR2_X1 U393 ( .A(n474), .B(n713), .Z(n354) );
  AND2_X2 U394 ( .A1(n387), .A2(n363), .ZN(n541) );
  XNOR2_X2 U395 ( .A(n577), .B(n501), .ZN(n639) );
  XNOR2_X2 U396 ( .A(n500), .B(G469), .ZN(n577) );
  NOR2_X1 U397 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X2 U398 ( .A1(n653), .A2(n652), .ZN(n413) );
  INV_X1 U399 ( .A(n398), .ZN(n377) );
  INV_X2 U400 ( .A(G116), .ZN(n443) );
  AND2_X1 U401 ( .A1(n553), .A2(n412), .ZN(n618) );
  XNOR2_X1 U402 ( .A(n416), .B(KEYINPUT42), .ZN(n731) );
  INV_X1 U403 ( .A(KEYINPUT16), .ZN(n531) );
  XNOR2_X1 U404 ( .A(n439), .B(n414), .ZN(n729) );
  XNOR2_X1 U405 ( .A(n413), .B(n574), .ZN(n666) );
  INV_X1 U406 ( .A(n564), .ZN(n634) );
  XNOR2_X1 U407 ( .A(n475), .B(n476), .ZN(n518) );
  XNOR2_X1 U408 ( .A(n483), .B(n482), .ZN(n533) );
  XOR2_X1 U409 ( .A(G137), .B(G140), .Z(n492) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(G119), .ZN(n444) );
  XNOR2_X1 U411 ( .A(G113), .B(G101), .ZN(n487) );
  INV_X1 U412 ( .A(KEYINPUT82), .ZN(n426) );
  XNOR2_X1 U413 ( .A(n381), .B(n557), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n381), .B(n557), .ZN(n672) );
  NAND2_X2 U415 ( .A1(n404), .A2(n625), .ZN(n572) );
  XNOR2_X2 U416 ( .A(n456), .B(n364), .ZN(n404) );
  AND2_X1 U417 ( .A1(n411), .A2(n586), .ZN(n457) );
  AND2_X1 U418 ( .A1(n650), .A2(n458), .ZN(n411) );
  XNOR2_X1 U419 ( .A(n384), .B(KEYINPUT73), .ZN(n676) );
  NOR2_X2 U420 ( .A1(n728), .A2(n618), .ZN(n383) );
  INV_X2 U421 ( .A(n590), .ZN(n597) );
  XNOR2_X1 U422 ( .A(n490), .B(n489), .ZN(n637) );
  NOR2_X1 U423 ( .A1(G902), .A2(n609), .ZN(n490) );
  XNOR2_X1 U424 ( .A(n533), .B(n463), .ZN(n491) );
  XNOR2_X1 U425 ( .A(n464), .B(G134), .ZN(n463) );
  INV_X1 U426 ( .A(G131), .ZN(n464) );
  XNOR2_X1 U427 ( .A(n451), .B(G953), .ZN(n717) );
  XNOR2_X1 U428 ( .A(n454), .B(n354), .ZN(n696) );
  XNOR2_X1 U429 ( .A(n455), .B(n477), .ZN(n454) );
  XNOR2_X1 U430 ( .A(n512), .B(n511), .ZN(n689) );
  XNOR2_X1 U431 ( .A(n510), .B(n466), .ZN(n511) );
  XNOR2_X1 U432 ( .A(n491), .B(n492), .ZN(n712) );
  INV_X1 U433 ( .A(KEYINPUT22), .ZN(n388) );
  NOR2_X1 U434 ( .A1(n628), .A2(n613), .ZN(n402) );
  XNOR2_X1 U435 ( .A(n391), .B(n390), .ZN(n389) );
  INV_X1 U436 ( .A(KEYINPUT44), .ZN(n390) );
  XNOR2_X1 U437 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n453) );
  NAND2_X1 U438 ( .A1(n518), .A2(G221), .ZN(n455) );
  XNOR2_X1 U439 ( .A(n375), .B(n528), .ZN(n374) );
  XNOR2_X1 U440 ( .A(KEYINPUT103), .B(n567), .ZN(n568) );
  AND2_X1 U441 ( .A1(n377), .A2(n625), .ZN(n394) );
  INV_X1 U442 ( .A(KEYINPUT0), .ZN(n419) );
  INV_X1 U443 ( .A(KEYINPUT91), .ZN(n452) );
  XNOR2_X1 U444 ( .A(n480), .B(n360), .ZN(n564) );
  XNOR2_X1 U445 ( .A(n430), .B(n491), .ZN(n609) );
  BUF_X1 U446 ( .A(n717), .Z(n418) );
  INV_X1 U447 ( .A(n696), .ZN(n449) );
  XNOR2_X1 U448 ( .A(n437), .B(n519), .ZN(n694) );
  XNOR2_X1 U449 ( .A(n521), .B(n520), .ZN(n437) );
  XNOR2_X1 U450 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U451 ( .A(n499), .B(n495), .ZN(n427) );
  NOR2_X1 U452 ( .A1(n674), .A2(n673), .ZN(n675) );
  INV_X1 U453 ( .A(KEYINPUT80), .ZN(n423) );
  INV_X1 U454 ( .A(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U455 ( .A(n434), .B(KEYINPUT97), .ZN(n654) );
  OR2_X1 U456 ( .A1(n629), .A2(n625), .ZN(n434) );
  XNOR2_X1 U457 ( .A(n515), .B(KEYINPUT4), .ZN(n483) );
  XNOR2_X1 U458 ( .A(G128), .B(G119), .ZN(n472) );
  XOR2_X1 U459 ( .A(KEYINPUT24), .B(G110), .Z(n473) );
  XNOR2_X1 U460 ( .A(n442), .B(G104), .ZN(n530) );
  INV_X1 U461 ( .A(G122), .ZN(n442) );
  XNOR2_X1 U462 ( .A(G140), .B(G143), .ZN(n504) );
  XOR2_X1 U463 ( .A(KEYINPUT94), .B(G131), .Z(n505) );
  XNOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n508) );
  XOR2_X1 U465 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n509) );
  XNOR2_X1 U466 ( .A(n525), .B(n527), .ZN(n375) );
  XNOR2_X1 U467 ( .A(n526), .B(n428), .ZN(n527) );
  XNOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n428) );
  NAND2_X1 U469 ( .A1(n634), .A2(n633), .ZN(n638) );
  XNOR2_X1 U470 ( .A(n436), .B(G478), .ZN(n544) );
  OR2_X1 U471 ( .A1(n694), .A2(G902), .ZN(n436) );
  XNOR2_X1 U472 ( .A(G146), .B(G137), .ZN(n484) );
  INV_X1 U473 ( .A(KEYINPUT81), .ZN(n600) );
  INV_X1 U474 ( .A(G953), .ZN(n704) );
  XOR2_X1 U475 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n476) );
  XOR2_X1 U476 ( .A(G101), .B(G107), .Z(n497) );
  XNOR2_X1 U477 ( .A(G146), .B(G104), .ZN(n494) );
  NAND2_X1 U478 ( .A1(G237), .A2(G234), .ZN(n538) );
  AND2_X1 U479 ( .A1(n568), .A2(n625), .ZN(n591) );
  OR2_X1 U480 ( .A1(n637), .A2(n415), .ZN(n563) );
  NAND2_X1 U481 ( .A1(n404), .A2(n629), .ZN(n631) );
  XNOR2_X1 U482 ( .A(n397), .B(KEYINPUT109), .ZN(n724) );
  AND2_X1 U483 ( .A1(n568), .A2(n394), .ZN(n569) );
  XNOR2_X1 U484 ( .A(n438), .B(KEYINPUT83), .ZN(n414) );
  INV_X1 U485 ( .A(KEYINPUT35), .ZN(n438) );
  XNOR2_X1 U486 ( .A(n435), .B(KEYINPUT96), .ZN(n629) );
  NOR2_X1 U487 ( .A1(n545), .A2(n546), .ZN(n435) );
  NOR2_X1 U488 ( .A1(n576), .A2(n634), .ZN(n412) );
  NOR2_X1 U489 ( .A1(n550), .A2(n403), .ZN(n613) );
  NAND2_X1 U490 ( .A1(n459), .A2(n637), .ZN(n403) );
  NAND2_X1 U491 ( .A1(n553), .A2(n421), .ZN(n554) );
  XNOR2_X1 U492 ( .A(n401), .B(n367), .ZN(n400) );
  INV_X1 U493 ( .A(KEYINPUT122), .ZN(n445) );
  XNOR2_X1 U494 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U495 ( .A(n693), .B(n694), .ZN(n385) );
  INV_X1 U496 ( .A(KEYINPUT60), .ZN(n460) );
  XNOR2_X1 U497 ( .A(n686), .B(n687), .ZN(n382) );
  INV_X1 U498 ( .A(KEYINPUT56), .ZN(n408) );
  XNOR2_X1 U499 ( .A(n424), .B(n423), .ZN(n677) );
  XNOR2_X1 U500 ( .A(n637), .B(n366), .ZN(n566) );
  INV_X1 U501 ( .A(n566), .ZN(n421) );
  AND2_X1 U502 ( .A1(n396), .A2(n622), .ZN(n356) );
  XNOR2_X1 U503 ( .A(KEYINPUT14), .B(n538), .ZN(n357) );
  XNOR2_X1 U504 ( .A(G902), .B(KEYINPUT15), .ZN(n358) );
  XOR2_X1 U505 ( .A(n380), .B(n379), .Z(n359) );
  XOR2_X1 U506 ( .A(n479), .B(n481), .Z(n360) );
  AND2_X1 U507 ( .A1(n507), .A2(G214), .ZN(n361) );
  AND2_X1 U508 ( .A1(n586), .A2(n458), .ZN(n362) );
  AND2_X1 U509 ( .A1(n469), .A2(n421), .ZN(n363) );
  XOR2_X1 U510 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n364) );
  AND2_X1 U511 ( .A1(n537), .A2(n357), .ZN(n365) );
  XOR2_X1 U512 ( .A(KEYINPUT99), .B(KEYINPUT6), .Z(n366) );
  INV_X1 U513 ( .A(n585), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n418), .A2(G952), .ZN(n697) );
  INV_X1 U515 ( .A(n697), .ZN(n447) );
  XOR2_X1 U516 ( .A(n609), .B(n468), .Z(n367) );
  XNOR2_X1 U517 ( .A(n712), .B(n427), .ZN(n682) );
  XOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT84), .Z(n368) );
  XNOR2_X1 U519 ( .A(n691), .B(n690), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n376), .A2(n447), .ZN(n409) );
  XNOR2_X1 U521 ( .A(n410), .B(n681), .ZN(n376) );
  NAND2_X1 U522 ( .A1(n650), .A2(n649), .ZN(n653) );
  INV_X1 U523 ( .A(n649), .ZN(n415) );
  XNOR2_X2 U524 ( .A(n369), .B(n532), .ZN(n699) );
  XNOR2_X2 U525 ( .A(n370), .B(n530), .ZN(n369) );
  XNOR2_X2 U526 ( .A(n529), .B(n531), .ZN(n370) );
  XNOR2_X1 U527 ( .A(n487), .B(KEYINPUT3), .ZN(n371) );
  NAND2_X1 U528 ( .A1(n372), .A2(n539), .ZN(n540) );
  NAND2_X1 U529 ( .A1(n372), .A2(n645), .ZN(n548) );
  XNOR2_X1 U530 ( .A(n372), .B(KEYINPUT89), .ZN(n550) );
  XNOR2_X2 U531 ( .A(n420), .B(n419), .ZN(n372) );
  NAND2_X1 U532 ( .A1(n359), .A2(n356), .ZN(n378) );
  NAND2_X1 U533 ( .A1(n654), .A2(KEYINPUT47), .ZN(n380) );
  NAND2_X1 U534 ( .A1(n590), .A2(n649), .ZN(n398) );
  NAND2_X1 U535 ( .A1(n462), .A2(n447), .ZN(n461) );
  NAND2_X1 U536 ( .A1(n400), .A2(n447), .ZN(n399) );
  NAND2_X1 U537 ( .A1(n448), .A2(n447), .ZN(n446) );
  XOR2_X1 U538 ( .A(KEYINPUT5), .B(n425), .Z(n485) );
  XNOR2_X1 U539 ( .A(n486), .B(n488), .ZN(n395) );
  XNOR2_X1 U540 ( .A(n395), .B(n532), .ZN(n430) );
  NAND2_X1 U541 ( .A1(n584), .A2(n583), .ZN(n396) );
  NOR2_X2 U542 ( .A1(n582), .A2(n581), .ZN(n623) );
  XNOR2_X1 U543 ( .A(n407), .B(n368), .ZN(n405) );
  NOR2_X1 U544 ( .A1(n378), .A2(n724), .ZN(n406) );
  XNOR2_X2 U545 ( .A(n541), .B(KEYINPUT32), .ZN(n728) );
  NAND2_X1 U546 ( .A1(n389), .A2(n556), .ZN(n381) );
  NOR2_X1 U547 ( .A1(n382), .A2(n697), .ZN(G54) );
  XNOR2_X1 U548 ( .A(n383), .B(KEYINPUT86), .ZN(n393) );
  NOR2_X2 U549 ( .A1(n672), .A2(n607), .ZN(n384) );
  NOR2_X1 U550 ( .A1(n385), .A2(n697), .ZN(G63) );
  XNOR2_X1 U551 ( .A(n386), .B(KEYINPUT34), .ZN(n441) );
  NAND2_X1 U552 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U553 ( .A(n729), .ZN(n392) );
  NAND2_X1 U554 ( .A1(n570), .A2(n593), .ZN(n397) );
  XNOR2_X2 U555 ( .A(n398), .B(KEYINPUT19), .ZN(n580) );
  XNOR2_X1 U556 ( .A(n399), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U557 ( .A1(n695), .A2(G472), .ZN(n401) );
  XNOR2_X1 U558 ( .A(n402), .B(KEYINPUT92), .ZN(n551) );
  NAND2_X1 U559 ( .A1(n405), .A2(n406), .ZN(n433) );
  NAND2_X1 U560 ( .A1(n731), .A2(n730), .ZN(n407) );
  XNOR2_X1 U561 ( .A(n409), .B(n408), .ZN(G51) );
  NAND2_X1 U562 ( .A1(n695), .A2(G210), .ZN(n410) );
  XNOR2_X2 U563 ( .A(n572), .B(n571), .ZN(n730) );
  NOR2_X1 U564 ( .A1(n551), .A2(n654), .ZN(n552) );
  NAND2_X1 U565 ( .A1(n457), .A2(n459), .ZN(n456) );
  XNOR2_X2 U566 ( .A(n597), .B(KEYINPUT38), .ZN(n650) );
  XNOR2_X1 U567 ( .A(n417), .B(KEYINPUT28), .ZN(n579) );
  AND2_X1 U568 ( .A1(n575), .A2(n576), .ZN(n417) );
  NAND2_X1 U569 ( .A1(n564), .A2(n633), .ZN(n565) );
  NAND2_X1 U570 ( .A1(n599), .A2(n631), .ZN(n422) );
  NAND2_X1 U571 ( .A1(n675), .A2(n676), .ZN(n424) );
  XNOR2_X1 U572 ( .A(n606), .B(n426), .ZN(n607) );
  XNOR2_X1 U573 ( .A(n461), .B(n460), .ZN(G60) );
  NOR2_X1 U574 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U575 ( .A1(n431), .A2(n632), .ZN(n605) );
  XNOR2_X1 U576 ( .A(n433), .B(n432), .ZN(n431) );
  INV_X1 U577 ( .A(KEYINPUT48), .ZN(n432) );
  NAND2_X1 U578 ( .A1(n441), .A2(n440), .ZN(n439) );
  INV_X1 U579 ( .A(n587), .ZN(n440) );
  XNOR2_X2 U580 ( .A(n443), .B(G107), .ZN(n529) );
  XNOR2_X1 U581 ( .A(n446), .B(n445), .ZN(G66) );
  NAND2_X1 U582 ( .A1(n695), .A2(G217), .ZN(n450) );
  INV_X1 U583 ( .A(KEYINPUT64), .ZN(n451) );
  NAND2_X1 U584 ( .A1(n459), .A2(n362), .ZN(n588) );
  XNOR2_X1 U585 ( .A(n549), .B(n452), .ZN(n459) );
  BUF_X1 U586 ( .A(n695), .Z(n692) );
  INV_X1 U587 ( .A(n577), .ZN(n578) );
  AND2_X1 U588 ( .A1(G210), .A2(n536), .ZN(n465) );
  XOR2_X1 U589 ( .A(n509), .B(n508), .Z(n466) );
  XOR2_X1 U590 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n467) );
  XNOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n468) );
  NOR2_X1 U592 ( .A1(n639), .A2(n634), .ZN(n469) );
  XNOR2_X1 U593 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n522), .B(KEYINPUT100), .ZN(n573) );
  INV_X1 U595 ( .A(n533), .ZN(n534) );
  INV_X1 U596 ( .A(n573), .ZN(n652) );
  XNOR2_X1 U597 ( .A(n680), .B(n467), .ZN(n681) );
  XOR2_X1 U598 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n471) );
  XNOR2_X1 U599 ( .A(KEYINPUT74), .B(KEYINPUT90), .ZN(n470) );
  XNOR2_X1 U600 ( .A(n471), .B(n470), .ZN(n481) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n492), .Z(n477) );
  NAND2_X1 U603 ( .A1(G234), .A2(n717), .ZN(n475) );
  NOR2_X1 U604 ( .A1(n696), .A2(G902), .ZN(n480) );
  NAND2_X1 U605 ( .A1(G234), .A2(n358), .ZN(n478) );
  XNOR2_X1 U606 ( .A(KEYINPUT20), .B(n478), .ZN(n502) );
  NAND2_X1 U607 ( .A1(G217), .A2(n502), .ZN(n479) );
  XOR2_X2 U608 ( .A(G128), .B(G143), .Z(n515) );
  XOR2_X1 U609 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n482) );
  XNOR2_X1 U610 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U611 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U612 ( .A1(n507), .A2(G210), .ZN(n488) );
  XNOR2_X1 U613 ( .A(KEYINPUT72), .B(G472), .ZN(n489) );
  INV_X1 U614 ( .A(KEYINPUT76), .ZN(n493) );
  NAND2_X1 U615 ( .A1(G227), .A2(n717), .ZN(n496) );
  XOR2_X1 U616 ( .A(n497), .B(n496), .Z(n498) );
  XOR2_X1 U617 ( .A(G110), .B(KEYINPUT88), .Z(n698) );
  XNOR2_X1 U618 ( .A(KEYINPUT71), .B(n698), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n498), .B(n525), .ZN(n499) );
  NOR2_X1 U620 ( .A1(n682), .A2(G902), .ZN(n500) );
  XNOR2_X1 U621 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n501) );
  INV_X1 U622 ( .A(n639), .ZN(n593) );
  NAND2_X1 U623 ( .A1(n502), .A2(G221), .ZN(n503) );
  XOR2_X1 U624 ( .A(KEYINPUT21), .B(n503), .Z(n633) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .ZN(n514) );
  XNOR2_X1 U626 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U627 ( .A(n530), .B(G113), .ZN(n510) );
  NOR2_X1 U628 ( .A1(G902), .A2(n689), .ZN(n513) );
  XOR2_X1 U629 ( .A(KEYINPUT7), .B(G134), .Z(n517) );
  XNOR2_X1 U630 ( .A(n529), .B(n515), .ZN(n516) );
  XNOR2_X1 U631 ( .A(n517), .B(n516), .ZN(n521) );
  XOR2_X1 U632 ( .A(G122), .B(KEYINPUT9), .Z(n520) );
  NAND2_X1 U633 ( .A1(G217), .A2(n518), .ZN(n519) );
  NAND2_X1 U634 ( .A1(n633), .A2(n573), .ZN(n523) );
  XNOR2_X1 U635 ( .A(n523), .B(KEYINPUT101), .ZN(n539) );
  NOR2_X1 U636 ( .A1(G898), .A2(n704), .ZN(n701) );
  NAND2_X1 U637 ( .A1(n701), .A2(G902), .ZN(n524) );
  NAND2_X1 U638 ( .A1(G952), .A2(n704), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n524), .A2(n559), .ZN(n537) );
  NAND2_X1 U640 ( .A1(G224), .A2(n418), .ZN(n528) );
  NAND2_X1 U641 ( .A1(n680), .A2(n358), .ZN(n535) );
  OR2_X1 U642 ( .A1(G902), .A2(G237), .ZN(n536) );
  XNOR2_X2 U643 ( .A(n535), .B(n465), .ZN(n590) );
  NAND2_X1 U644 ( .A1(G214), .A2(n536), .ZN(n649) );
  NAND2_X1 U645 ( .A1(n546), .A2(n544), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n547), .A2(n566), .ZN(n543) );
  XOR2_X1 U647 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n542) );
  XNOR2_X1 U648 ( .A(n543), .B(n542), .ZN(n665) );
  INV_X1 U649 ( .A(n544), .ZN(n545) );
  AND2_X1 U650 ( .A1(n546), .A2(n545), .ZN(n625) );
  INV_X1 U651 ( .A(n637), .ZN(n576) );
  AND2_X1 U652 ( .A1(n547), .A2(n576), .ZN(n645) );
  XNOR2_X1 U653 ( .A(KEYINPUT31), .B(n548), .ZN(n628) );
  NOR2_X1 U654 ( .A1(n577), .A2(n638), .ZN(n549) );
  XNOR2_X1 U655 ( .A(KEYINPUT98), .B(n552), .ZN(n555) );
  NOR2_X1 U656 ( .A1(n564), .A2(n554), .ZN(n610) );
  NOR2_X1 U657 ( .A1(n555), .A2(n610), .ZN(n556) );
  INV_X1 U658 ( .A(KEYINPUT45), .ZN(n557) );
  NOR2_X1 U659 ( .A1(n418), .A2(G900), .ZN(n558) );
  NAND2_X1 U660 ( .A1(G902), .A2(n558), .ZN(n560) );
  NAND2_X1 U661 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U662 ( .A1(n357), .A2(n561), .ZN(n585) );
  XOR2_X1 U663 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n562) );
  XNOR2_X1 U664 ( .A(n563), .B(n562), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n585), .A2(n565), .ZN(n575) );
  NAND2_X1 U666 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U667 ( .A(KEYINPUT36), .B(n569), .ZN(n570) );
  XOR2_X1 U668 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n571) );
  XNOR2_X1 U669 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n574) );
  NAND2_X1 U670 ( .A1(n579), .A2(n578), .ZN(n582) );
  INV_X1 U671 ( .A(n580), .ZN(n581) );
  XOR2_X1 U672 ( .A(n623), .B(KEYINPUT47), .Z(n584) );
  NAND2_X1 U673 ( .A1(n623), .A2(n654), .ZN(n583) );
  NOR2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n622) );
  XNOR2_X1 U676 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n591), .A2(n649), .ZN(n592) );
  NOR2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT105), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n598), .A2(n597), .ZN(n632) );
  INV_X1 U682 ( .A(n605), .ZN(n599) );
  NOR2_X1 U683 ( .A1(KEYINPUT2), .A2(n601), .ZN(n602) );
  NOR2_X1 U684 ( .A1(n602), .A2(n358), .ZN(n608) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(n631), .ZN(n603) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n603), .Z(n604) );
  AND2_X2 U687 ( .A1(n608), .A2(n676), .ZN(n695) );
  XOR2_X1 U688 ( .A(G101), .B(n610), .Z(G3) );
  XOR2_X1 U689 ( .A(G104), .B(KEYINPUT111), .Z(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n625), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n612), .B(n611), .ZN(G6) );
  XNOR2_X1 U692 ( .A(G107), .B(KEYINPUT112), .ZN(n617) );
  XOR2_X1 U693 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n615) );
  NAND2_X1 U694 ( .A1(n613), .A2(n629), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(G9) );
  XOR2_X1 U697 ( .A(n618), .B(G110), .Z(G12) );
  XOR2_X1 U698 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n620) );
  NAND2_X1 U699 ( .A1(n623), .A2(n629), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(n621) );
  XOR2_X1 U701 ( .A(G128), .B(n621), .Z(G30) );
  XNOR2_X1 U702 ( .A(G143), .B(n622), .ZN(G45) );
  NAND2_X1 U703 ( .A1(n623), .A2(n625), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(G146), .ZN(G48) );
  NAND2_X1 U705 ( .A1(n628), .A2(n625), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT114), .ZN(n627) );
  XNOR2_X1 U707 ( .A(G113), .B(n627), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(n425), .ZN(G18) );
  XNOR2_X1 U710 ( .A(G134), .B(n631), .ZN(G36) );
  XNOR2_X1 U711 ( .A(G140), .B(n632), .ZN(G42) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n635), .B(KEYINPUT49), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n642) );
  AND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT50), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT116), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT51), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT117), .B(n647), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n666), .A2(n648), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U727 ( .A1(n665), .A2(n657), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT52), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT118), .ZN(n663) );
  NAND2_X1 U731 ( .A1(G952), .A2(n357), .ZN(n662) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U733 ( .A1(G953), .A2(n664), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT119), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n678) );
  INV_X1 U737 ( .A(KEYINPUT2), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n670), .A2(n716), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n671), .B(KEYINPUT79), .ZN(n674) );
  INV_X1 U740 ( .A(n355), .ZN(n703) );
  NOR2_X1 U741 ( .A1(KEYINPUT2), .A2(n703), .ZN(n673) );
  XNOR2_X1 U742 ( .A(KEYINPUT53), .B(n679), .ZN(G75) );
  XOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n684) );
  XNOR2_X1 U744 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U746 ( .A(n682), .B(n685), .Z(n687) );
  NAND2_X1 U747 ( .A1(n692), .A2(G469), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n695), .A2(G475), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT59), .B(KEYINPUT87), .Z(n688) );
  NAND2_X1 U750 ( .A1(G478), .A2(n692), .ZN(n693) );
  XOR2_X1 U751 ( .A(n699), .B(n698), .Z(n700) );
  XNOR2_X1 U752 ( .A(KEYINPUT123), .B(n700), .ZN(n702) );
  NOR2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n711) );
  NAND2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n705) );
  XNOR2_X1 U756 ( .A(KEYINPUT61), .B(n705), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n706), .A2(G898), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U759 ( .A(n709), .B(KEYINPUT124), .ZN(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(G69) );
  XOR2_X1 U761 ( .A(n713), .B(n712), .Z(n719) );
  INV_X1 U762 ( .A(n719), .ZN(n714) );
  XNOR2_X1 U763 ( .A(KEYINPUT125), .B(n714), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n718), .A2(n418), .ZN(n723) );
  XNOR2_X1 U766 ( .A(G227), .B(n719), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(G900), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n721), .A2(G953), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n723), .A2(n722), .ZN(G72) );
  XOR2_X1 U770 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n726) );
  XNOR2_X1 U771 ( .A(n724), .B(G125), .ZN(n725) );
  XNOR2_X1 U772 ( .A(n726), .B(n725), .ZN(G27) );
  XOR2_X1 U773 ( .A(G119), .B(KEYINPUT126), .Z(n727) );
  XNOR2_X1 U774 ( .A(n728), .B(n727), .ZN(G21) );
  XOR2_X1 U775 ( .A(n729), .B(G122), .Z(G24) );
  XNOR2_X1 U776 ( .A(n730), .B(G131), .ZN(G33) );
  XNOR2_X1 U777 ( .A(n731), .B(G137), .ZN(G39) );
endmodule

