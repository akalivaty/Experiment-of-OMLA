//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT82), .A2(G101), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT82), .A2(G101), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n200), .A2(new_n191), .A3(new_n194), .A4(new_n195), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT0), .A3(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n213));
  NAND3_X1  g027(.A1(new_n196), .A2(G101), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n203), .A2(new_n216), .A3(G128), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n207), .B(G146), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n208), .B2(new_n210), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G104), .B(G107), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT84), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n190), .A2(G107), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n193), .A2(G104), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n228), .B(G101), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n224), .A2(new_n232), .A3(KEYINPUT10), .A4(new_n201), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n215), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n217), .A2(new_n223), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n232), .A3(new_n201), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT10), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT85), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n234), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT64), .B(new_n244), .C1(new_n245), .C2(G137), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G134), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT64), .B1(new_n249), .B2(new_n244), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(new_n245), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n248), .A2(G134), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(G131), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(G137), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n246), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT88), .B1(new_n243), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n215), .A2(new_n233), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n227), .A2(new_n231), .B1(new_n273), .B2(new_n200), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n274), .C2(new_n236), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n241), .B1(new_n237), .B2(new_n238), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT88), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n269), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n272), .B(new_n270), .C1(new_n275), .C2(new_n276), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n240), .A2(new_n242), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT86), .A3(new_n270), .A4(new_n272), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT81), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(KEYINPUT89), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT89), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n271), .A2(new_n279), .B1(new_n283), .B2(new_n285), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n292), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n293), .B1(new_n283), .B2(new_n285), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n237), .B1(new_n224), .B2(new_n274), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT87), .A3(new_n269), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT12), .Z(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n294), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G469), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n292), .B1(new_n301), .B2(new_n286), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n280), .B2(new_n298), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n309), .B2(G469), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n189), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G237), .ZN(new_n315));
  INV_X1    g129(.A(G237), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n317));
  OAI211_X1 g131(.A(G214), .B(new_n288), .C1(new_n315), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n207), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(G237), .ZN(new_n321));
  AOI21_X1  g135(.A(G953), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n313), .B1(new_n324), .B2(G131), .ZN(new_n325));
  AOI211_X1 g139(.A(KEYINPUT96), .B(new_n267), .C1(new_n319), .C2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT17), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT98), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n209), .ZN(new_n338));
  OAI211_X1 g152(.A(G146), .B(new_n332), .C1(new_n336), .C2(new_n330), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT75), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n341), .A3(new_n209), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n325), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT17), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n324), .A2(new_n313), .A3(G131), .ZN(new_n346));
  INV_X1    g160(.A(new_n324), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n267), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT98), .B(KEYINPUT17), .C1(new_n325), .C2(new_n326), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n329), .A2(new_n343), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT18), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n352), .B2(new_n267), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n324), .A2(KEYINPUT18), .A3(G131), .ZN(new_n354));
  INV_X1    g168(.A(new_n336), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n209), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n336), .B2(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n209), .B2(new_n355), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G113), .B(G122), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT97), .B(G104), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n351), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n336), .B(KEYINPUT19), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n339), .B1(new_n367), .B2(G146), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n325), .A2(new_n326), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n348), .ZN(new_n370));
  INV_X1    g184(.A(new_n361), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n312), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  AOI211_X1 g190(.A(KEYINPUT20), .B(new_n376), .C1(new_n366), .C2(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n351), .A2(new_n361), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n364), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n379), .B2(new_n366), .ZN(new_n380));
  INV_X1    g194(.A(G475), .ZN(new_n381));
  OAI22_X1  g195(.A1(new_n375), .A2(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  INV_X1    g197(.A(G122), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n384), .A2(KEYINPUT99), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(KEYINPUT99), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(KEYINPUT67), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n390), .A3(G122), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n387), .A2(new_n392), .A3(G107), .ZN(new_n393));
  XNOR2_X1  g207(.A(G128), .B(G143), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n245), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n387), .B1(new_n391), .B2(KEYINPUT14), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n193), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G107), .B1(new_n387), .B2(new_n392), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT13), .B1(new_n222), .B2(G143), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(new_n245), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n403), .A2(new_n394), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n394), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n393), .A2(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n187), .A2(new_n407), .A3(G953), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n400), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT100), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n400), .B2(new_n406), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT100), .B(new_n409), .C1(new_n400), .C2(new_n406), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n305), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n382), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n311), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(G234), .A2(G237), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(G952), .A3(new_n288), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(G902), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n388), .A2(new_n390), .A3(G119), .ZN(new_n428));
  INV_X1    g242(.A(G119), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G116), .ZN(new_n430));
  INV_X1    g244(.A(G113), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT2), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT2), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G113), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT68), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n428), .A2(new_n435), .A3(new_n438), .A4(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n428), .A2(KEYINPUT5), .A3(new_n430), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n431), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n274), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(new_n430), .ZN(new_n447));
  INV_X1    g261(.A(new_n435), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n437), .A2(new_n439), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n202), .A2(new_n214), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n445), .B(new_n446), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n204), .A2(new_n211), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G125), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n217), .A2(new_n221), .A3(new_n334), .A4(new_n223), .ZN(new_n454));
  INV_X1    g268(.A(G224), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G953), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n453), .B2(new_n454), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n446), .B(KEYINPUT8), .Z(new_n463));
  AOI22_X1  g277(.A1(new_n437), .A2(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(new_n274), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(new_n445), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n305), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT93), .B(new_n305), .C1(new_n462), .C2(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  INV_X1    g286(.A(new_n450), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n447), .A2(new_n448), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n440), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n473), .A2(new_n475), .B1(new_n464), .B2(new_n274), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n472), .B1(new_n476), .B2(new_n446), .ZN(new_n477));
  INV_X1    g291(.A(new_n446), .ZN(new_n478));
  INV_X1    g292(.A(new_n445), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n449), .A2(new_n450), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT90), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n481), .A4(new_n451), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT91), .B(KEYINPUT6), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n478), .B(new_n483), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n453), .A2(new_n454), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n456), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n482), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n471), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT94), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G214), .B1(G237), .B2(G902), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n471), .A2(new_n489), .A3(new_n492), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT95), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n494), .A2(new_n499), .A3(new_n495), .A4(new_n496), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n427), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n420), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n452), .B1(new_n260), .B2(new_n268), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n249), .B1(new_n261), .B2(G134), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G131), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n268), .A2(new_n224), .A3(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n503), .A2(new_n506), .A3(KEYINPUT30), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n262), .A2(new_n266), .A3(new_n267), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n267), .B1(new_n262), .B2(new_n266), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n212), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n268), .A2(new_n224), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n475), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n449), .A3(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n322), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n475), .B1(new_n503), .B2(new_n506), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(new_n524), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n521), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT30), .B1(new_n503), .B2(new_n506), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n449), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n516), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(new_n521), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT71), .B1(new_n535), .B2(new_n515), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n514), .A2(new_n516), .A3(new_n522), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT31), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n530), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT32), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n523), .A2(new_n529), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n535), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n538), .B1(new_n537), .B2(KEYINPUT31), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n541), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n525), .A2(new_n516), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n527), .A3(new_n522), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n305), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n514), .A2(new_n516), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n556), .B2(new_n521), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(KEYINPUT72), .A3(new_n527), .A4(new_n522), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n305), .C1(new_n552), .C2(new_n553), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n543), .A2(new_n549), .B1(G472), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n407), .B1(G234), .B2(new_n305), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(G119), .B(G128), .Z(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT74), .B1(new_n429), .B2(G128), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n576), .A2(KEYINPUT23), .B1(new_n429), .B2(G128), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT23), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT74), .B(new_n578), .C1(new_n429), .C2(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(G110), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n340), .A2(new_n342), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT78), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n573), .A2(new_n574), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n580), .B2(G110), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n339), .A3(new_n359), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n583), .B1(new_n582), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n572), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  INV_X1    g405(.A(new_n572), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n568), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n305), .A3(new_n593), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT79), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n566), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n600), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n589), .A2(KEYINPUT25), .A3(new_n593), .A4(new_n305), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(KEYINPUT79), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n597), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n565), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n502), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n200), .B(KEYINPUT101), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT102), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n610), .B(new_n612), .ZN(G3));
  NAND2_X1  g427(.A1(new_n306), .A2(new_n310), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n540), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n547), .A2(new_n541), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n614), .A2(new_n617), .A3(new_n607), .A4(new_n188), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n311), .A2(KEYINPUT103), .A3(new_n607), .A4(new_n617), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n413), .A2(new_n622), .A3(new_n414), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n410), .A2(KEYINPUT33), .A3(new_n412), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(G478), .A3(new_n305), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n415), .A2(new_n416), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n373), .A2(new_n374), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT20), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n373), .A2(new_n312), .A3(new_n374), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n366), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n365), .B1(new_n351), .B2(new_n361), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n305), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G475), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n628), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n427), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n494), .A2(new_n638), .A3(new_n495), .A4(new_n496), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n382), .A2(new_n627), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT104), .B1(new_n643), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n620), .A2(new_n621), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  OAI211_X1 g462(.A(new_n636), .B(new_n418), .C1(new_n375), .C2(new_n377), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n639), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n620), .A2(new_n621), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n590), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n567), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n604), .A2(KEYINPUT79), .A3(new_n605), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n602), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n617), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n502), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n658), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n543), .A2(new_n549), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n564), .A2(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n497), .ZN(new_n667));
  INV_X1    g481(.A(new_n418), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n422), .B(KEYINPUT105), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n425), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n382), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n666), .A2(new_n667), .A3(new_n311), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(new_n672), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n311), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  INV_X1    g493(.A(G472), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n550), .B2(new_n521), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n537), .A2(new_n681), .B1(G472), .B2(G902), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n664), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n494), .A2(new_n496), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT107), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n382), .A2(new_n418), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n663), .A2(new_n495), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n678), .A2(new_n679), .A3(new_n684), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n672), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n382), .A2(new_n627), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n666), .A2(new_n667), .A3(new_n311), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  AND3_X1   g512(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n189), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n641), .B1(new_n637), .B2(new_n640), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n643), .A2(KEYINPUT104), .A3(new_n639), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n609), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n701), .A2(new_n609), .A3(new_n650), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NOR4_X1   g522(.A1(new_n699), .A2(new_n700), .A3(new_n497), .A4(new_n189), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n632), .A2(new_n668), .A3(new_n636), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n565), .A2(new_n710), .A3(new_n663), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n711), .A3(new_n638), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND2_X1  g527(.A1(new_n303), .A2(new_n305), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n188), .A3(new_n306), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n535), .A2(new_n515), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n541), .B1(new_n717), .B2(new_n530), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n607), .A2(new_n615), .A3(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n716), .A2(new_n427), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n630), .A2(new_n631), .B1(G475), .B2(new_n635), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n668), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n382), .A2(KEYINPUT109), .A3(new_n418), .ZN(new_n724));
  AND4_X1   g538(.A1(KEYINPUT110), .A2(new_n723), .A3(new_n667), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n497), .B1(new_n689), .B2(new_n721), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n720), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND3_X1  g543(.A1(new_n615), .A2(new_n658), .A3(new_n718), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n695), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n701), .A2(new_n667), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT111), .B(G125), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G27));
  XOR2_X1   g548(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n735));
  NAND2_X1  g549(.A1(new_n311), .A2(new_n696), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n548), .B1(new_n547), .B2(new_n541), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n542), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n665), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n495), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n494), .B2(new_n496), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n607), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n735), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n741), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n565), .A2(new_n746), .A3(new_n608), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n311), .A4(new_n696), .ZN(new_n748));
  OAI211_X1 g562(.A(KEYINPUT113), .B(new_n735), .C1(new_n736), .C2(new_n742), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  AND3_X1   g565(.A1(new_n673), .A2(new_n614), .A3(new_n188), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n747), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n311), .A2(new_n673), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n742), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NOR2_X1   g572(.A1(new_n382), .A2(new_n628), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT43), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n617), .A2(new_n663), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT44), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n746), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n298), .A2(new_n280), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n301), .A2(new_n286), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(new_n292), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n304), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n309), .A2(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n307), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n306), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n188), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n760), .A2(KEYINPUT44), .A3(new_n761), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n763), .A2(new_n774), .A3(new_n676), .A4(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT115), .B(G137), .Z(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G39));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  OAI221_X1 g593(.A(new_n188), .B1(KEYINPUT116), .B2(new_n779), .C1(new_n771), .C2(new_n772), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n739), .A2(new_n695), .A3(new_n746), .A4(new_n607), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT116), .B(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n781), .C1(new_n774), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(new_n699), .A2(new_n700), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT49), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n495), .A2(new_n688), .A3(new_n188), .A4(new_n759), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n684), .A2(new_n608), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n760), .A2(new_n670), .ZN(new_n790));
  INV_X1    g604(.A(new_n719), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n701), .A2(new_n740), .A3(new_n688), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT117), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n796), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n794), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n716), .A2(new_n746), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n423), .A3(new_n788), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n722), .A3(new_n628), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n801), .A2(new_n760), .A3(new_n670), .ZN(new_n804));
  INV_X1    g618(.A(new_n730), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n785), .A2(new_n189), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n782), .B1(new_n773), .B2(new_n188), .ZN(new_n809));
  INV_X1    g623(.A(new_n780), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n760), .A2(new_n670), .A3(new_n791), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n746), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n797), .A2(new_n800), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n709), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT119), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(KEYINPUT119), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n804), .A2(new_n609), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT48), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n288), .A2(G952), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n802), .B2(new_n637), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT120), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n803), .A2(new_n806), .A3(KEYINPUT51), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n798), .B2(new_n794), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n811), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n813), .B1(new_n811), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n822), .A2(new_n824), .A3(new_n835), .A4(new_n826), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n817), .A2(new_n828), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n427), .B(new_n643), .C1(new_n498), .C2(new_n500), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n620), .A2(new_n838), .A3(new_n621), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n427), .B(new_n649), .C1(new_n498), .C2(new_n500), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n620), .A2(new_n621), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n420), .B(new_n501), .C1(new_n609), .C2(new_n659), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n658), .A2(new_n672), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n311), .A2(new_n684), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n723), .A2(new_n667), .A3(new_n724), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n726), .A2(KEYINPUT110), .A3(new_n724), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n732), .A2(new_n674), .A3(new_n697), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n732), .A2(new_n674), .A3(new_n697), .ZN(new_n853));
  INV_X1    g667(.A(new_n845), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n725), .B2(new_n727), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n843), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n749), .A2(new_n748), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n609), .A2(new_n311), .A3(new_n696), .A4(new_n741), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT113), .B1(new_n860), .B2(new_n735), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n609), .B(new_n701), .C1(new_n645), .C2(new_n650), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n728), .A2(new_n712), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n311), .A2(new_n741), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n565), .A2(new_n710), .A3(new_n663), .A4(new_n672), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n731), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n755), .A2(new_n742), .A3(new_n754), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT114), .B1(new_n752), .B2(new_n747), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n862), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n732), .A2(new_n674), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(KEYINPUT52), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n843), .A2(new_n852), .A3(new_n857), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n712), .A2(new_n704), .A3(new_n707), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n739), .A2(new_n419), .A3(new_n658), .A4(new_n694), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n695), .B2(new_n730), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n753), .A2(new_n756), .B1(new_n879), .B2(new_n865), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n750), .A2(new_n728), .A3(new_n877), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n872), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n873), .A2(KEYINPUT52), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n872), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n858), .A2(new_n871), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n888), .B2(new_n883), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n837), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n789), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n288), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n305), .B1(new_n875), .B2(new_n882), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(new_n492), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n488), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n895), .A2(new_n492), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n902), .A4(new_n899), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(G51));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n307), .ZN(new_n909));
  INV_X1    g723(.A(new_n884), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n883), .B1(new_n875), .B2(new_n882), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n303), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n768), .A2(new_n769), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT123), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n895), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n893), .B1(new_n913), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n895), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n373), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT124), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G60));
  NOR2_X1   g738(.A1(new_n910), .A2(new_n911), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n623), .A2(new_n624), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n894), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n889), .A2(new_n928), .B1(new_n623), .B2(new_n624), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n407), .A2(new_n305), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n875), .B2(new_n882), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n655), .B(KEYINPUT126), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n595), .A2(new_n596), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n894), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n933), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n938), .A2(new_n943), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n894), .A4(new_n940), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G66));
  NAND3_X1  g762(.A1(new_n843), .A2(new_n728), .A3(new_n877), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(G953), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n426), .B2(new_n455), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n897), .B1(G898), .B2(new_n288), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  NOR2_X1   g772(.A1(new_n507), .A2(new_n513), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n367), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n671), .B2(new_n288), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n609), .B1(new_n725), .B2(new_n727), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n774), .A2(new_n676), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n783), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n776), .A2(new_n757), .A3(new_n853), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n862), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(new_n288), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n692), .A2(new_n853), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n677), .B1(new_n643), .B2(new_n649), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n747), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n970), .A2(new_n776), .A3(new_n783), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n960), .B1(new_n973), .B2(new_n288), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n967), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n967), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT63), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n521), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n973), .B2(new_n949), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n556), .B(new_n522), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n522), .A2(new_n980), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n966), .B2(new_n950), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n894), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n888), .A2(new_n983), .A3(new_n980), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G57));
endmodule


