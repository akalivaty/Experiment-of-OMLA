

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XOR2_X2 U326 ( .A(KEYINPUT38), .B(n448), .Z(n499) );
  XOR2_X1 U327 ( .A(n426), .B(n345), .Z(n518) );
  XOR2_X1 U328 ( .A(G8GAT), .B(G78GAT), .Z(n294) );
  XNOR2_X1 U329 ( .A(n403), .B(n294), .ZN(n409) );
  XNOR2_X1 U330 ( .A(n337), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U331 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U332 ( .A(n339), .B(n338), .ZN(n340) );
  NOR2_X1 U333 ( .A1(n468), .A2(n492), .ZN(n575) );
  XNOR2_X1 U334 ( .A(n465), .B(KEYINPUT48), .ZN(n549) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n475) );
  XNOR2_X1 U336 ( .A(n475), .B(KEYINPUT58), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n449), .B(G43GAT), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n477), .B(n476), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT82), .B(G71GAT), .Z(n296) );
  XNOR2_X1 U341 ( .A(KEYINPUT65), .B(KEYINPUT84), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U343 ( .A(G176GAT), .B(KEYINPUT81), .Z(n298) );
  XNOR2_X1 U344 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n300), .B(n299), .Z(n311) );
  INV_X1 U347 ( .A(KEYINPUT19), .ZN(n301) );
  NAND2_X1 U348 ( .A1(n301), .A2(KEYINPUT17), .ZN(n304) );
  INV_X1 U349 ( .A(KEYINPUT17), .ZN(n302) );
  NAND2_X1 U350 ( .A1(n302), .A2(KEYINPUT19), .ZN(n303) );
  NAND2_X1 U351 ( .A1(n304), .A2(n303), .ZN(n306) );
  XNOR2_X1 U352 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n339) );
  XOR2_X1 U354 ( .A(G99GAT), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n339), .B(n309), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U359 ( .A(G127GAT), .B(KEYINPUT20), .Z(n313) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U362 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U363 ( .A(KEYINPUT80), .B(G134GAT), .Z(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(n318), .ZN(n359) );
  XOR2_X1 U367 ( .A(G169GAT), .B(n359), .Z(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n531) );
  INV_X1 U369 ( .A(n531), .ZN(n473) );
  XOR2_X1 U370 ( .A(G29GAT), .B(KEYINPUT7), .Z(n322) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G36GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U373 ( .A(G50GAT), .B(KEYINPUT8), .Z(n323) );
  XOR2_X1 U374 ( .A(n324), .B(n323), .Z(n446) );
  XOR2_X1 U375 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n326) );
  XNOR2_X1 U376 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(n327), .ZN(n331) );
  XOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .Z(n427) );
  XOR2_X1 U380 ( .A(n427), .B(G92GAT), .Z(n329) );
  NAND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(G218GAT), .B(G162GAT), .Z(n370) );
  XOR2_X1 U385 ( .A(n332), .B(n370), .Z(n334) );
  XNOR2_X1 U386 ( .A(G134GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n446), .B(n335), .ZN(n560) );
  XOR2_X1 U389 ( .A(n560), .B(KEYINPUT36), .Z(n588) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n336), .B(G64GAT), .ZN(n426) );
  XOR2_X1 U392 ( .A(G169GAT), .B(G8GAT), .Z(n439) );
  XOR2_X1 U393 ( .A(G197GAT), .B(KEYINPUT21), .Z(n369) );
  XNOR2_X1 U394 ( .A(n439), .B(n369), .ZN(n344) );
  XOR2_X1 U395 ( .A(G183GAT), .B(G211GAT), .Z(n400) );
  AND2_X1 U396 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U397 ( .A(n400), .B(n340), .Z(n342) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U401 ( .A(KEYINPUT27), .B(n518), .Z(n388) );
  XOR2_X1 U402 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n347) );
  XNOR2_X1 U403 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U405 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n349) );
  XNOR2_X1 U406 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n374) );
  XOR2_X1 U408 ( .A(n374), .B(KEYINPUT89), .Z(n351) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n358) );
  XOR2_X1 U411 ( .A(G57GAT), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(G148GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(G127GAT), .B(G155GAT), .Z(n399) );
  XOR2_X1 U415 ( .A(n354), .B(n399), .Z(n356) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(G85GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n516) );
  INV_X1 U421 ( .A(n516), .ZN(n492) );
  NAND2_X1 U422 ( .A1(n388), .A2(n492), .ZN(n363) );
  XOR2_X1 U423 ( .A(KEYINPUT90), .B(n363), .Z(n548) );
  XOR2_X1 U424 ( .A(G148GAT), .B(G106GAT), .Z(n365) );
  XNOR2_X1 U425 ( .A(G204GAT), .B(G78GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U427 ( .A(KEYINPUT73), .B(n366), .Z(n435) );
  XOR2_X1 U428 ( .A(G155GAT), .B(G211GAT), .Z(n368) );
  XNOR2_X1 U429 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U431 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n372) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U434 ( .A(n373), .B(KEYINPUT87), .Z(n380) );
  INV_X1 U435 ( .A(G22GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n377) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n378), .B(G50GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U441 ( .A(n382), .B(n381), .Z(n383) );
  XOR2_X1 U442 ( .A(n435), .B(n383), .Z(n469) );
  XOR2_X1 U443 ( .A(n469), .B(KEYINPUT28), .Z(n498) );
  INV_X1 U444 ( .A(n498), .ZN(n527) );
  NAND2_X1 U445 ( .A1(n548), .A2(n527), .ZN(n530) );
  XNOR2_X1 U446 ( .A(n530), .B(KEYINPUT91), .ZN(n384) );
  NAND2_X1 U447 ( .A1(n384), .A2(n531), .ZN(n396) );
  INV_X1 U448 ( .A(KEYINPUT26), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n473), .A2(n469), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(KEYINPUT92), .B(n387), .Z(n576) );
  AND2_X1 U452 ( .A1(n388), .A2(n576), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n389), .B(KEYINPUT93), .ZN(n393) );
  INV_X1 U454 ( .A(n518), .ZN(n495) );
  NAND2_X1 U455 ( .A1(n473), .A2(n495), .ZN(n390) );
  NAND2_X1 U456 ( .A1(n469), .A2(n390), .ZN(n391) );
  XOR2_X1 U457 ( .A(KEYINPUT25), .B(n391), .Z(n392) );
  NAND2_X1 U458 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U459 ( .A1(n394), .A2(n516), .ZN(n395) );
  NAND2_X1 U460 ( .A1(n396), .A2(n395), .ZN(n481) );
  XOR2_X1 U461 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n398) );
  XNOR2_X1 U462 ( .A(KEYINPUT12), .B(KEYINPUT78), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n411) );
  XOR2_X1 U464 ( .A(KEYINPUT15), .B(n399), .Z(n402) );
  XNOR2_X1 U465 ( .A(G64GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U467 ( .A(G1GAT), .B(KEYINPUT67), .Z(n405) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(G15GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n442) );
  XNOR2_X1 U470 ( .A(n442), .B(KEYINPUT79), .ZN(n407) );
  AND2_X1 U471 ( .A1(G231GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n411), .B(n410), .Z(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT70), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U475 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U477 ( .A(KEYINPUT69), .B(n414), .Z(n431) );
  XNOR2_X1 U478 ( .A(n415), .B(n431), .ZN(n457) );
  NAND2_X1 U479 ( .A1(n481), .A2(n457), .ZN(n416) );
  XNOR2_X1 U480 ( .A(KEYINPUT96), .B(n416), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n588), .A2(n417), .ZN(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT37), .B(KEYINPUT97), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n515) );
  XOR2_X1 U484 ( .A(KEYINPUT75), .B(KEYINPUT71), .Z(n421) );
  XNOR2_X1 U485 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U487 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n423) );
  XNOR2_X1 U488 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U490 ( .A(n425), .B(n424), .Z(n433) );
  XOR2_X1 U491 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U492 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n582) );
  XOR2_X1 U497 ( .A(KEYINPUT66), .B(G113GAT), .Z(n437) );
  XNOR2_X1 U498 ( .A(G141GAT), .B(G197GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U504 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n578) );
  XOR2_X1 U507 ( .A(n578), .B(KEYINPUT68), .Z(n564) );
  NOR2_X1 U508 ( .A1(n582), .A2(n564), .ZN(n482) );
  NAND2_X1 U509 ( .A1(n515), .A2(n482), .ZN(n448) );
  NAND2_X1 U510 ( .A1(n473), .A2(n499), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n449) );
  INV_X1 U512 ( .A(n560), .ZN(n542) );
  XOR2_X1 U513 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n471) );
  XOR2_X1 U514 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n467) );
  XOR2_X1 U515 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n452) );
  XNOR2_X1 U516 ( .A(n452), .B(n582), .ZN(n554) );
  NAND2_X1 U517 ( .A1(n578), .A2(n554), .ZN(n453) );
  XNOR2_X1 U518 ( .A(KEYINPUT46), .B(n453), .ZN(n454) );
  INV_X1 U519 ( .A(n457), .ZN(n478) );
  XOR2_X1 U520 ( .A(KEYINPUT110), .B(n478), .Z(n573) );
  NAND2_X1 U521 ( .A1(n454), .A2(n573), .ZN(n455) );
  NOR2_X1 U522 ( .A1(n560), .A2(n455), .ZN(n456) );
  XNOR2_X1 U523 ( .A(KEYINPUT47), .B(n456), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n588), .A2(n457), .ZN(n458) );
  XNOR2_X1 U525 ( .A(n458), .B(KEYINPUT45), .ZN(n460) );
  INV_X1 U526 ( .A(n582), .ZN(n459) );
  NAND2_X1 U527 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U528 ( .A(n461), .B(KEYINPUT111), .ZN(n462) );
  NAND2_X1 U529 ( .A1(n462), .A2(n564), .ZN(n463) );
  NAND2_X1 U530 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U531 ( .A1(n549), .A2(n495), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U533 ( .A1(n575), .A2(n469), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n472), .B(KEYINPUT55), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n474), .A2(n473), .ZN(n572) );
  NOR2_X1 U537 ( .A1(n542), .A2(n572), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n542), .A2(n478), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  AND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n502) );
  NAND2_X1 U541 ( .A1(n482), .A2(n502), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n516), .A2(n490), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U545 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U546 ( .A1(n518), .A2(n490), .ZN(n486) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n531), .A2(n490), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT95), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NOR2_X1 U552 ( .A1(n527), .A2(n490), .ZN(n491) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U555 ( .A1(n492), .A2(n499), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT98), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT100), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n554), .ZN(n566) );
  NOR2_X1 U564 ( .A1(n566), .A2(n578), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n514), .A2(n502), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT102), .B(n503), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n516), .A2(n510), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n518), .A2(n510), .ZN(n508) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n510), .A2(n531), .ZN(n509) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n527), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n516), .A2(n526), .ZN(n517) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n531), .A2(n526), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n525) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(n529), .B(n528), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n549), .A2(n532), .ZN(n543) );
  NOR2_X1 U597 ( .A1(n564), .A2(n543), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n566), .A2(n543), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n573), .A2(n543), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n545) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U615 ( .A(n576), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT118), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n578), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U621 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n478), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n572), .ZN(n565) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n572), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .ZN(n589) );
  INV_X1 U643 ( .A(n589), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n582), .A2(n585), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n478), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

