//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  OR3_X1    g004(.A1(new_n190), .A2(KEYINPUT16), .A3(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G146), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G146), .B1(new_n189), .B2(new_n191), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n201), .C1(G119), .C2(new_n200), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  AOI22_X1  g018(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n192), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n189), .A2(KEYINPUT74), .A3(G146), .A4(new_n191), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n188), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n202), .A2(G110), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n204), .A2(KEYINPUT72), .A3(new_n203), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT72), .B1(new_n204), .B2(new_n203), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT73), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT73), .A4(new_n216), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n223), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n207), .B2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n230), .B2(G902), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT25), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G234), .B2(new_n232), .ZN(new_n236));
  INV_X1    g050(.A(new_n230), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(G902), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n234), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G472), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n211), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G134), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n259), .B2(KEYINPUT11), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n255), .B2(G134), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(G137), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n259), .A2(KEYINPUT11), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n254), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n250), .A2(KEYINPUT1), .A3(new_n200), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n273));
  AOI21_X1  g087(.A(G128), .B1(new_n247), .B2(new_n249), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n275), .A2(new_n211), .A3(G143), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n211), .A2(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(KEYINPUT68), .C1(new_n244), .C2(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n272), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n255), .A2(KEYINPUT67), .A3(G134), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n258), .B2(G137), .ZN(new_n284));
  OAI211_X1 g098(.A(G131), .B(new_n282), .C1(new_n284), .C2(new_n256), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n265), .A2(new_n285), .ZN(new_n286));
  OAI22_X1  g100(.A1(new_n270), .A2(new_n271), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n265), .ZN(new_n288));
  INV_X1    g102(.A(new_n254), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(new_n271), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n242), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G116), .B(G119), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT2), .B(G113), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT69), .B1(new_n269), .B2(new_n265), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n244), .A2(new_n275), .A3(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n248), .A2(G146), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n200), .B1(new_n300), .B2(new_n278), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT68), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n274), .A2(new_n273), .A3(new_n276), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n265), .A3(new_n285), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n291), .A2(new_n295), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n298), .A2(new_n294), .A3(new_n305), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n294), .A4(new_n305), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT27), .Z(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G101), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n314), .B(new_n315), .Z(new_n316));
  NAND4_X1  g130(.A1(new_n307), .A2(new_n310), .A3(new_n311), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT31), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n310), .A2(new_n311), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n316), .A4(new_n307), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n308), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT28), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n295), .B1(new_n287), .B2(new_n290), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n310), .A2(new_n325), .A3(new_n311), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n316), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n241), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n316), .ZN(new_n331));
  AND4_X1   g145(.A1(new_n310), .A2(new_n307), .A3(new_n311), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g147(.A(G902), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n335));
  INV_X1    g149(.A(new_n324), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n316), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n298), .A2(new_n305), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n310), .B(new_n311), .C1(new_n294), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT28), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n341), .B2(new_n336), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n334), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n330), .A2(KEYINPUT32), .B1(new_n343), .B2(G472), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n329), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n318), .B(new_n321), .C1(new_n327), .C2(new_n316), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n241), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n240), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT9), .B(G234), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n232), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G221), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT76), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n277), .A2(new_n280), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n299), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n361));
  AOI21_X1  g175(.A(G101), .B1(new_n360), .B2(G107), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G104), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n360), .A2(G107), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n367), .A2(new_n369), .B1(G101), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n299), .A2(new_n301), .A3(new_n279), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(G101), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n359), .A2(new_n373), .B1(new_n377), .B2(new_n357), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n361), .A2(new_n365), .A3(new_n371), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G101), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n379), .A2(KEYINPUT79), .A3(new_n380), .A4(G101), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n254), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n380), .B1(new_n379), .B2(G101), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n374), .A2(KEYINPUT78), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT78), .B1(new_n374), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n296), .A2(new_n297), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n377), .B1(new_n304), .B2(new_n373), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n288), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT12), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G140), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n224), .A2(G227), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n297), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT12), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n392), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n391), .A2(new_n394), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n393), .A2(KEYINPUT12), .B1(new_n401), .B2(new_n392), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(KEYINPUT80), .A3(new_n391), .A4(new_n398), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n378), .A2(new_n389), .ZN(new_n409));
  INV_X1    g223(.A(new_n390), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n391), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT81), .B1(new_n412), .B2(new_n397), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n378), .A2(new_n389), .A3(new_n390), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n390), .B1(new_n378), .B2(new_n389), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT81), .B(new_n397), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n408), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n232), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n397), .B1(new_n414), .B2(new_n415), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n416), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n425), .B2(new_n408), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n419), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n412), .A2(new_n398), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n406), .A2(new_n391), .A3(new_n397), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n232), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G469), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n356), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(G475), .A2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n312), .A2(G214), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n248), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n312), .B(G214), .C1(KEYINPUT84), .C2(G143), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT18), .A2(G131), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n188), .A2(new_n211), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n441), .A2(new_n442), .B1(new_n212), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n440), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n445), .A2(KEYINPUT85), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT85), .B1(new_n445), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n439), .A2(new_n261), .A3(new_n440), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n261), .B1(new_n439), .B2(new_n440), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(G131), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n261), .A3(new_n440), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n458), .A2(KEYINPUT19), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(KEYINPUT19), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n188), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n188), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n209), .B(new_n210), .C1(G146), .C2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n449), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(G113), .B(G122), .Z(new_n465));
  XOR2_X1   g279(.A(KEYINPUT88), .B(G104), .Z(new_n466));
  XOR2_X1   g280(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n470), .A3(new_n455), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n452), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT89), .B1(new_n452), .B2(KEYINPUT17), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n195), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n467), .A3(new_n449), .ZN(new_n475));
  AOI211_X1 g289(.A(KEYINPUT20), .B(new_n436), .C1(new_n469), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n475), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n435), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n478), .B2(new_n435), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n475), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n467), .B1(new_n474), .B2(new_n449), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n232), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT92), .B1(new_n200), .B2(G143), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n248), .A3(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n200), .A2(G143), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n494), .A2(new_n258), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(G116), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G116), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(KEYINPUT91), .A3(G122), .ZN(new_n501));
  OAI22_X1  g315(.A1(new_n499), .A2(new_n501), .B1(G116), .B2(new_n498), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n502), .A2(G107), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(G107), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n495), .B1(new_n494), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n494), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT93), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n494), .A2(new_n510), .A3(new_n506), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n505), .B1(new_n258), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n505), .B(KEYINPUT94), .C1(new_n258), .C2(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n499), .A2(new_n501), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n504), .B1(KEYINPUT14), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n258), .B1(new_n494), .B2(new_n495), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n364), .A2(KEYINPUT14), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n496), .A2(new_n520), .B1(new_n502), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n353), .A2(G217), .A3(new_n224), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n526), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n517), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n232), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n528), .B1(new_n517), .B2(new_n524), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n523), .B(new_n526), .C1(new_n515), .C2(new_n516), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n232), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G952), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G953), .ZN(new_n541));
  NAND2_X1  g355(.A1(G234), .A2(G237), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(G902), .A3(G953), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n490), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G214), .B1(G237), .B2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n294), .B1(new_n383), .B2(new_n384), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n387), .B2(new_n388), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n500), .A2(KEYINPUT5), .A3(G119), .ZN(new_n554));
  INV_X1    g368(.A(G113), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n293), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n553), .A2(new_n556), .B1(new_n557), .B2(new_n292), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n373), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G122), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n552), .A2(new_n561), .A3(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n254), .A2(G125), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n304), .B2(G125), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n571), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT7), .B1(new_n568), .B2(G953), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n561), .B(KEYINPUT8), .ZN(new_n576));
  INV_X1    g390(.A(new_n559), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n373), .A2(new_n558), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n567), .A2(new_n574), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n581), .B2(new_n564), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G210), .B1(G237), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT83), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n583), .B(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n549), .A2(new_n550), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n351), .A2(new_n434), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n348), .A2(new_n232), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(new_n346), .A3(new_n349), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n433), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n421), .B2(new_n428), .ZN(new_n597));
  NOR4_X1   g411(.A1(new_n595), .A2(new_n240), .A3(new_n597), .A4(new_n356), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n573), .A2(new_n582), .A3(KEYINPUT95), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n585), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n550), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT95), .B1(new_n573), .B2(new_n582), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n584), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n531), .A2(new_n232), .ZN(new_n607));
  INV_X1    g421(.A(new_n537), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(new_n531), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n530), .A2(KEYINPUT33), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT33), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(G478), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n490), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n606), .A2(new_n613), .A3(new_n548), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  AOI22_X1  g431(.A1(new_n484), .A2(new_n480), .B1(G475), .B2(new_n488), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n548), .B(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n539), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  AND2_X1   g438(.A1(new_n346), .A2(new_n349), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n234), .A2(new_n236), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n222), .B(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n238), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n625), .A2(KEYINPUT98), .A3(new_n593), .A4(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n593), .A2(new_n632), .A3(new_n346), .A4(new_n349), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n633), .A2(new_n636), .A3(new_n434), .A4(new_n589), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT99), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n546), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n543), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n489), .B(new_n643), .C1(new_n483), .C2(new_n476), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n534), .B2(new_n538), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n602), .A2(new_n645), .A3(new_n605), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n630), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n238), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n344), .A2(new_n350), .B1(new_n626), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n648), .A2(new_n651), .A3(new_n434), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(new_n643), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n434), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n319), .A2(new_n307), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n316), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n232), .C1(new_n316), .C2(new_n340), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n330), .A2(KEYINPUT32), .B1(G472), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n350), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n588), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n490), .A2(new_n539), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n664), .A2(new_n603), .A3(new_n632), .A4(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n656), .A2(new_n657), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT102), .B(G143), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G45));
  INV_X1    g483(.A(new_n643), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n606), .A2(new_n613), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n651), .A2(new_n434), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI22_X1  g487(.A1(new_n424), .A2(new_n416), .B1(new_n405), .B2(new_n407), .ZN(new_n674));
  OAI21_X1  g488(.A(G469), .B1(new_n674), .B2(G902), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n427), .B1(new_n426), .B2(new_n419), .ZN(new_n676));
  NOR4_X1   g490(.A1(new_n674), .A2(KEYINPUT82), .A3(G469), .A4(G902), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n355), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n351), .A2(new_n614), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NAND3_X1  g496(.A1(new_n351), .A2(new_n621), .A3(new_n679), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  NOR2_X1   g498(.A1(new_n678), .A2(new_n606), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n651), .A2(new_n685), .A3(new_n549), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  NOR2_X1   g501(.A1(new_n606), .A2(new_n665), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n316), .B1(new_n341), .B2(new_n336), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n241), .B1(new_n322), .B2(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n593), .A2(new_n239), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n679), .A2(new_n688), .A3(new_n619), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT103), .B(G122), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G24));
  AND4_X1   g508(.A1(new_n490), .A2(new_n609), .A3(new_n612), .A4(new_n643), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n593), .A2(new_n632), .A3(new_n690), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n685), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G125), .ZN(G27));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n355), .B1(new_n597), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n701), .B(new_n433), .C1(new_n676), .C2(new_n677), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT105), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n433), .B1(new_n676), .B2(new_n677), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n706), .A2(KEYINPUT104), .B1(G221), .B2(new_n354), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n703), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n588), .A2(new_n603), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n343), .A2(G472), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n347), .B2(new_n329), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n239), .B(new_n695), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n705), .A2(new_n709), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  INV_X1    g531(.A(new_n710), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n355), .A3(new_n703), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n718), .B1(new_n720), .B2(KEYINPUT105), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n351), .A3(new_n709), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n261), .ZN(G33));
  NAND4_X1  g539(.A1(new_n721), .A2(new_n351), .A3(new_n645), .A4(new_n709), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  INV_X1    g541(.A(new_n490), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n612), .A3(new_n609), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n729), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n595), .A3(new_n632), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n430), .A2(new_n431), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n419), .B1(new_n739), .B2(KEYINPUT45), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(KEYINPUT45), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT46), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n429), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n355), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n747), .A2(new_n654), .A3(new_n710), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n736), .A2(new_n737), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n738), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(G137), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G39));
  NAND2_X1  g566(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n696), .A2(new_n718), .A3(new_n239), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n350), .A3(new_n344), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n643), .B(KEYINPUT112), .Z(new_n761));
  NOR2_X1   g575(.A1(new_n632), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n719), .A2(new_n355), .A3(new_n703), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT113), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n707), .A2(new_n765), .A3(new_n703), .A4(new_n762), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n662), .A2(new_n688), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n652), .A2(new_n672), .A3(new_n699), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n652), .A2(new_n672), .A3(new_n699), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n767), .A3(new_n766), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n717), .A3(new_n723), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n588), .A2(new_n550), .A3(new_n619), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n613), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n434), .A2(new_n239), .A3(new_n594), .A4(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n590), .A2(new_n778), .A3(KEYINPUT110), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT110), .B1(new_n590), .B2(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n539), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT111), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n728), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n776), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n434), .A2(new_n785), .A3(new_n239), .A4(new_n594), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n637), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n779), .A2(new_n780), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n705), .A2(new_n709), .A3(new_n698), .A4(new_n710), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n644), .B(new_n718), .C1(new_n783), .C2(new_n782), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n651), .A3(new_n434), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n680), .A2(new_n686), .A3(new_n683), .A4(new_n692), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n792), .A3(new_n726), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n760), .B1(new_n775), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n780), .A2(new_n787), .ZN(new_n796));
  INV_X1    g610(.A(new_n779), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n726), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n791), .A3(new_n789), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n724), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n652), .A2(new_n699), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n760), .B1(new_n803), .B2(KEYINPUT52), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n802), .A3(new_n774), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n795), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT53), .B1(new_n803), .B2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n800), .A2(new_n802), .A3(new_n774), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n806), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n774), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n724), .A3(new_n801), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n814), .B2(new_n800), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n775), .A2(new_n794), .A3(new_n808), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT54), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n795), .A2(new_n805), .A3(new_n806), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n735), .A2(new_n544), .A3(new_n691), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n718), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n756), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n356), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n429), .A2(new_n675), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n756), .A2(new_n823), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n735), .A2(new_n544), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n678), .A2(new_n718), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n662), .A2(new_n240), .A3(new_n543), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n609), .A2(new_n612), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n728), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n835), .A2(new_n697), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n679), .A2(new_n664), .A3(new_n603), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n841), .B1(new_n821), .B2(new_n842), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n821), .A2(new_n841), .A3(new_n842), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT51), .B1(new_n832), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n840), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n753), .A2(new_n755), .A3(new_n829), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n822), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n843), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .A4(KEYINPUT51), .ZN(new_n851));
  INV_X1    g665(.A(new_n685), .ZN(new_n852));
  OAI221_X1 g666(.A(new_n541), .B1(new_n613), .B2(new_n837), .C1(new_n821), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n713), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n240), .B1(new_n854), .B2(new_n344), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n833), .A2(new_n855), .A3(new_n834), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n846), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n812), .A2(new_n820), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n540), .A2(new_n224), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n729), .A2(new_n240), .A3(new_n356), .A4(new_n603), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT109), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT109), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n664), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OR4_X1    g686(.A1(new_n662), .A2(new_n869), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n864), .A2(KEYINPUT117), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n224), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n232), .B1(new_n795), .B2(new_n805), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n565), .A2(new_n572), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n570), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n885), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n742), .B(KEYINPUT57), .Z(new_n891));
  AOI21_X1  g705(.A(new_n806), .B1(new_n795), .B2(new_n805), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n807), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n418), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n881), .B(new_n740), .C1(KEYINPUT45), .C2(new_n739), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n879), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND2_X1  g710(.A1(KEYINPUT58), .A2(G475), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT119), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n881), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n478), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n899), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n880), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT120), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G60));
  NAND2_X1  g718(.A1(new_n610), .A2(new_n611), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n607), .B(KEYINPUT59), .Z(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n807), .C2(new_n892), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n880), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n812), .A2(new_n820), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n910), .B2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(G63));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n795), .A2(new_n805), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n235), .A2(new_n232), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n879), .B1(new_n919), .B2(new_n230), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n649), .A3(new_n918), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n913), .A2(KEYINPUT123), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(G66));
  OAI21_X1  g738(.A(G953), .B1(new_n547), .B2(new_n568), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n788), .A2(new_n793), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n883), .B1(G898), .B2(new_n224), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n747), .A2(new_n654), .A3(new_n688), .A4(new_n855), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n726), .A2(new_n750), .A3(new_n758), .A4(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n771), .B(KEYINPUT125), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n934), .A2(new_n717), .A3(new_n723), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n291), .A2(new_n306), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n462), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n641), .B2(new_n224), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n932), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n935), .A2(new_n667), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n718), .B1(new_n613), .B2(new_n784), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n351), .A3(new_n434), .A4(new_n654), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n750), .A2(new_n758), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n939), .B1(new_n948), .B2(new_n224), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT127), .Z(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n936), .B2(new_n927), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n879), .B1(new_n957), .B2(new_n332), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n948), .B2(new_n927), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n316), .A3(new_n658), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n795), .A2(new_n810), .ZN(new_n961));
  INV_X1    g775(.A(new_n332), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n659), .A4(new_n955), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n958), .A2(new_n960), .A3(new_n963), .ZN(G57));
endmodule


