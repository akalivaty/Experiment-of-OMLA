//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n205), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n220), .B(new_n225), .C1(G58), .C2(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n211), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n210), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n216), .B(new_n228), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n219), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT64), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT65), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n255), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n229), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n254), .A2(new_n256), .A3(new_n260), .A4(new_n229), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n209), .A2(G20), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n258), .A2(KEYINPUT71), .A3(new_n259), .A4(new_n261), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n264), .A2(G50), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n259), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n202), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n258), .A2(new_n261), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n203), .A2(G20), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n210), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n271), .B1(new_n272), .B2(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n267), .A2(new_n269), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n267), .A2(KEYINPUT9), .A3(new_n269), .A4(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT75), .ZN(new_n284));
  XOR2_X1   g0084(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT66), .B(G45), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n209), .B1(new_n286), .B2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  AND2_X1   g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n229), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n209), .C1(new_n286), .C2(G41), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n288), .A2(G274), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G226), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT3), .B(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G222), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G223), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n305), .B1(new_n246), .B2(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n290), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n294), .A2(KEYINPUT68), .A3(new_n299), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G200), .B2(new_n311), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n284), .A2(KEYINPUT77), .A3(new_n285), .A4(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n283), .A2(KEYINPUT75), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT75), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n281), .B2(new_n282), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n314), .B(new_n285), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT77), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n281), .A3(new_n282), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n315), .A2(new_n321), .B1(KEYINPUT10), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n311), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(new_n279), .C1(G169), .C2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n276), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT73), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G20), .B2(G77), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n331), .B1(new_n275), .B2(new_n274), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n270), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n268), .A2(new_n246), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n258), .A2(new_n261), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G77), .A3(new_n265), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n298), .A2(G244), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n294), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n303), .A2(G232), .A3(new_n304), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G107), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n342), .B(new_n346), .C1(new_n306), .C2(new_n223), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n345), .A2(new_n304), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G238), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(new_n342), .A3(KEYINPUT72), .A4(new_n346), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n352), .A3(new_n290), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT74), .B(new_n339), .C1(new_n354), .C2(G169), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT74), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n357));
  AOI21_X1  g0157(.A(G169), .B1(new_n341), .B2(new_n353), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n325), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n354), .A2(G190), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n357), .C1(new_n363), .C2(new_n354), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n323), .A2(new_n328), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n345), .B2(new_n210), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NOR4_X1   g0168(.A1(new_n343), .A2(new_n344), .A3(new_n368), .A4(G20), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n273), .A2(G159), .ZN(new_n371));
  AND2_X1   g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT81), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(G20), .C1(new_n372), .C2(new_n201), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n371), .A4(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n270), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n350), .A2(G226), .ZN(new_n383));
  NAND3_X1  g0183(.A1(KEYINPUT82), .A2(G33), .A3(G87), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n303), .A2(G223), .A3(new_n304), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT82), .ZN(new_n386));
  INV_X1    g0186(.A(G33), .ZN(new_n387));
  INV_X1    g0187(.A(G87), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n290), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n298), .A2(G232), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(G190), .A3(new_n294), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n275), .A2(new_n268), .ZN(new_n394));
  INV_X1    g0194(.A(new_n275), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n264), .A2(new_n265), .A3(new_n266), .A4(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n382), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n294), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G200), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OR3_X1    g0200(.A1(new_n397), .A2(new_n400), .A3(KEYINPUT17), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT17), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n382), .A2(new_n394), .A3(new_n396), .ZN(new_n404));
  INV_X1    g0204(.A(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n391), .A2(new_n325), .A3(new_n294), .A4(new_n392), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT83), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT18), .A4(new_n406), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n411), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(KEYINPUT80), .A2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n303), .A2(G226), .A3(new_n304), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n303), .A2(G232), .A3(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n387), .B2(new_n205), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G33), .A3(G97), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n290), .B1(new_n298), .B2(G238), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n294), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n424), .B2(new_n294), .ZN(new_n428));
  OAI211_X1 g0228(.A(G169), .B(new_n416), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G179), .A3(new_n426), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n405), .B1(new_n430), .B2(new_n426), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT80), .B(KEYINPUT14), .Z(new_n433));
  OAI211_X1 g0233(.A(new_n429), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n222), .A2(G20), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n435), .B1(new_n276), .B2(new_n246), .C1(new_n274), .C2(new_n202), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n270), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT11), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n337), .A2(G68), .A3(new_n265), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n435), .A2(G1), .A3(new_n212), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT12), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n434), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n427), .B2(new_n428), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n430), .A2(G190), .A3(new_n426), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n415), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n366), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n209), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n258), .A2(new_n259), .A3(new_n261), .A4(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n459));
  OAI21_X1  g0259(.A(G107), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n210), .A2(G107), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT23), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n388), .A2(KEYINPUT89), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n303), .A2(KEYINPUT22), .A3(new_n210), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n276), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G116), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n303), .A2(new_n210), .A3(new_n463), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(KEYINPUT24), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n462), .A3(new_n467), .A4(new_n464), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n474), .A3(new_n270), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n259), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT25), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n460), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n303), .A2(G250), .A3(new_n304), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n480), .C1(new_n306), .C2(new_n224), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n209), .B(G45), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n291), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n481), .A2(new_n290), .B1(new_n485), .B2(G264), .ZN(new_n486));
  INV_X1    g0286(.A(G274), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n484), .A2(new_n487), .A3(new_n290), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n486), .A2(new_n325), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(G169), .B1(new_n486), .B2(new_n489), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n478), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n218), .A2(G20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n257), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n210), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT84), .A2(G97), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT84), .A2(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n501), .B2(new_n387), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n494), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g0303(.A1(KEYINPUT84), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT84), .A2(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n210), .B(new_n497), .C1(new_n506), .C2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(KEYINPUT20), .A3(new_n257), .A4(new_n495), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n268), .A2(new_n218), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n509), .B(new_n510), .C1(new_n218), .C2(new_n457), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n303), .A2(G257), .A3(new_n304), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n345), .A2(G303), .ZN(new_n513));
  INV_X1    g0313(.A(G264), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n306), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n488), .B1(new_n515), .B2(new_n290), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n485), .A2(G270), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n405), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(KEYINPUT21), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT88), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n511), .A2(new_n518), .A3(new_n521), .A4(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n511), .B2(new_n518), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(G179), .A3(new_n517), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n526), .B2(new_n511), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n516), .A2(new_n517), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n312), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n511), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT86), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n207), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n504), .A2(KEYINPUT6), .A3(new_n206), .A4(new_n505), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT85), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n501), .A2(new_n544), .A3(KEYINPUT6), .A4(new_n206), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  OAI21_X1  g0347(.A(G107), .B1(new_n367), .B2(new_n369), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n273), .A2(G77), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n270), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n268), .A2(new_n205), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n458), .A2(new_n459), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n205), .ZN(new_n554));
  OAI211_X1 g0354(.A(G244), .B(new_n304), .C1(new_n343), .C2(new_n344), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n303), .A2(KEYINPUT4), .A3(G244), .A4(new_n304), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n303), .A2(G250), .A3(G1698), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n497), .A4(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n488), .B1(new_n560), .B2(new_n290), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n291), .A2(G257), .A3(new_n484), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n561), .A2(new_n325), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G169), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n554), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n312), .A3(new_n563), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n488), .B(new_n562), .C1(new_n560), .C2(new_n290), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(G200), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT87), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n337), .A2(new_n571), .A3(new_n259), .A4(new_n456), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G97), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n570), .A2(new_n575), .A3(new_n552), .A4(new_n551), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G238), .B(new_n304), .C1(new_n343), .C2(new_n344), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n343), .C2(new_n344), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n387), .C2(new_n218), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n290), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n209), .A2(G45), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n487), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(G250), .C1(new_n289), .C2(new_n229), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n325), .A2(new_n581), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n585), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n580), .B2(new_n290), .ZN(new_n588));
  AOI21_X1  g0388(.A(G169), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n329), .B1(new_n572), .B2(new_n573), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n501), .A2(G87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT19), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(new_n206), .B1(new_n593), .B2(new_n210), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n506), .B2(new_n276), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n303), .A2(new_n210), .A3(G68), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n270), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n329), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n259), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n590), .B1(new_n591), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n581), .A2(new_n312), .A3(new_n584), .A4(new_n585), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n583), .B(new_n587), .C1(new_n580), .C2(new_n290), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(G200), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n329), .A2(new_n268), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n553), .C2(new_n388), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n486), .A2(G190), .A3(new_n489), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n460), .A2(new_n475), .A3(new_n477), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n363), .B1(new_n486), .B2(new_n489), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n602), .B(new_n608), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n577), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n455), .A2(new_n493), .A3(new_n533), .A4(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n315), .A2(new_n321), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n322), .A2(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n450), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n447), .B1(new_n361), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n403), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n410), .A2(new_n412), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n328), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n493), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n478), .A2(new_n492), .A3(KEYINPUT90), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n523), .A3(new_n527), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n613), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT91), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n602), .A2(new_n554), .A3(new_n608), .A4(new_n566), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT93), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n630), .A2(new_n633), .A3(new_n631), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n602), .B(KEYINPUT92), .Z(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT91), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n627), .A2(new_n613), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n629), .A2(new_n636), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n623), .B1(new_n454), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT94), .ZN(G369));
  NOR2_X1   g0444(.A1(new_n212), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n209), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G343), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n511), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n533), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n523), .A2(new_n527), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n655), .A2(new_n652), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n610), .A2(new_n611), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n493), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n493), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n478), .A2(new_n652), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n493), .B2(new_n651), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n625), .A2(new_n626), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n651), .B(KEYINPUT95), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n660), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  NAND3_X1  g0472(.A1(new_n592), .A2(new_n206), .A3(new_n218), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n213), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n232), .B2(new_n676), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT96), .ZN(new_n680));
  INV_X1    g0480(.A(new_n493), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n528), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n602), .A2(new_n608), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n659), .A2(new_n683), .A3(new_n567), .A4(new_n576), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n613), .B(KEYINPUT96), .C1(new_n681), .C2(new_n528), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n630), .A2(new_n631), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n632), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n685), .A2(new_n686), .A3(new_n638), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT29), .A3(new_n651), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n627), .A2(new_n613), .A3(new_n639), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n639), .B1(new_n627), .B2(new_n613), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(KEYINPUT93), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n630), .A2(new_n633), .A3(new_n631), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n637), .B1(new_n696), .B2(new_n632), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n668), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n690), .B1(new_n698), .B2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n533), .A2(new_n613), .A3(new_n493), .A4(new_n669), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n604), .A2(new_n486), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n561), .A2(new_n563), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n525), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n486), .A2(new_n489), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(G179), .A3(new_n604), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n529), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n706), .A2(new_n707), .B1(new_n711), .B2(new_n529), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n651), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n701), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n700), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n679), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR2_X1   g0522(.A1(new_n213), .A2(new_n303), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n232), .B2(new_n286), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT98), .Z(new_n725));
  INV_X1    g0525(.A(new_n247), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n296), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n214), .A2(new_n303), .ZN(new_n728));
  XOR2_X1   g0528(.A(G355), .B(KEYINPUT97), .Z(new_n729));
  OAI221_X1 g0529(.A(new_n727), .B1(G116), .B2(new_n214), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n229), .B1(G20), .B2(new_n405), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT99), .Z(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(G20), .A2(G179), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n312), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n312), .A2(new_n363), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G322), .A2(new_n742), .B1(new_n745), .B2(G326), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n210), .A2(G179), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n312), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n312), .A3(new_n363), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n749), .A2(G283), .B1(new_n751), .B2(G329), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n740), .A2(new_n325), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n303), .B1(new_n754), .B2(G294), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n746), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n743), .A2(new_n747), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(G303), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n739), .A2(new_n312), .A3(new_n363), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n739), .A2(new_n312), .A3(G200), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI221_X1 g0563(.A(new_n759), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n744), .A2(new_n202), .ZN(new_n765));
  INV_X1    g0565(.A(G58), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n751), .A2(G159), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n741), .A2(new_n766), .B1(new_n767), .B2(KEYINPUT32), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(KEYINPUT32), .B2(new_n767), .ZN(new_n769));
  INV_X1    g0569(.A(new_n762), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G68), .B1(G97), .B2(new_n754), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n749), .A2(G107), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n303), .C1(new_n388), .C2(new_n757), .ZN(new_n773));
  INV_X1    g0573(.A(new_n761), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(G77), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n769), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n764), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n730), .A2(new_n737), .B1(new_n777), .B2(new_n734), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n209), .B1(new_n645), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n675), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n733), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n778), .B(new_n781), .C1(new_n656), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n657), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n656), .A2(G330), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(G396));
  NOR2_X1   g0587(.A1(new_n357), .A2(new_n651), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n361), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n361), .B2(new_n364), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n698), .B(new_n791), .Z(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(new_n720), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n720), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(new_n784), .A3(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G116), .A2(new_n774), .B1(new_n770), .B2(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n345), .B1(new_n757), .B2(new_n206), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n388), .A2(new_n748), .B1(new_n750), .B2(new_n760), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(G97), .C2(new_n754), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n742), .A2(G294), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n745), .A2(G303), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n796), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n762), .A2(new_n272), .B1(new_n744), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G159), .B2(new_n774), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n741), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n222), .A2(new_n748), .B1(new_n750), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n754), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n303), .B1(new_n811), .B2(new_n766), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(G50), .C2(new_n758), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n802), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n734), .A2(new_n731), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(new_n734), .B1(new_n246), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n781), .C1(new_n791), .C2(new_n732), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n795), .A2(new_n818), .ZN(G384));
  NAND3_X1  g0619(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n701), .A2(new_n820), .A3(new_n717), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n455), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT105), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n382), .A2(new_n396), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n824), .A2(new_n399), .A3(new_n393), .A4(new_n394), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n404), .A2(new_n650), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n408), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT104), .ZN(new_n829));
  INV_X1    g0629(.A(new_n397), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(new_n399), .B1(new_n404), .B2(new_n650), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT104), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n826), .A4(new_n408), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n382), .A2(new_n394), .A3(new_n396), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n649), .B1(new_n397), .B2(new_n400), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT37), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT103), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT103), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(KEYINPUT37), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n827), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n415), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  INV_X1    g0646(.A(new_n838), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n829), .B2(new_n833), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n827), .B1(new_n403), .B2(new_n621), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n446), .A2(new_n652), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n447), .A2(new_n450), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n446), .B(new_n652), .C1(new_n618), .C2(new_n434), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n791), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n821), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n851), .A2(new_n858), .A3(KEYINPUT40), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n829), .A2(new_n833), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n839), .A2(new_n841), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n844), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n846), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n857), .B1(new_n863), .B2(new_n845), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n859), .B1(new_n864), .B2(KEYINPUT40), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n823), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(G330), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n700), .A2(new_n455), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n623), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n447), .A2(new_n652), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n863), .B2(new_n845), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n845), .A2(new_n850), .A3(new_n871), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n410), .A2(new_n412), .A3(new_n649), .ZN(new_n875));
  INV_X1    g0675(.A(new_n855), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n641), .A2(new_n669), .A3(new_n791), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n361), .A2(new_n652), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n863), .A2(new_n845), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n869), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n867), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n209), .B2(new_n645), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n218), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n230), .C1(KEYINPUT35), .C2(new_n546), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n222), .B2(G50), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n202), .A2(KEYINPUT102), .A3(G68), .ZN(new_n892));
  OAI21_X1  g0692(.A(G77), .B1(new_n766), .B2(new_n222), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n891), .B(new_n892), .C1(new_n232), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n212), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT106), .Z(G367));
  OAI22_X1  g0697(.A1(new_n811), .A2(new_n222), .B1(new_n748), .B2(new_n246), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n345), .B(new_n898), .C1(G137), .C2(new_n751), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n758), .A2(G58), .ZN(new_n900));
  AOI22_X1  g0700(.A1(G50), .A2(new_n774), .B1(new_n770), .B2(G159), .ZN(new_n901));
  AOI22_X1  g0701(.A1(G143), .A2(new_n745), .B1(new_n742), .B2(G150), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n904));
  INV_X1    g0704(.A(G317), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n904), .B1(new_n905), .B2(new_n750), .C1(new_n506), .C2(new_n748), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n303), .B(new_n906), .C1(G311), .C2(new_n745), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT46), .B1(new_n758), .B2(G116), .ZN(new_n908));
  INV_X1    g0708(.A(G303), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n908), .A2(KEYINPUT109), .B1(new_n741), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(KEYINPUT109), .B2(new_n908), .ZN(new_n911));
  AOI22_X1  g0711(.A1(G283), .A2(new_n774), .B1(new_n770), .B2(G294), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n811), .A2(new_n206), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT47), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n784), .B1(new_n916), .B2(new_n734), .ZN(new_n917));
  INV_X1    g0717(.A(new_n723), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n737), .B1(new_n214), .B2(new_n329), .C1(new_n241), .C2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT108), .Z(new_n920));
  NAND2_X1  g0720(.A1(new_n574), .A2(G87), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n651), .B1(new_n921), .B2(new_n607), .ZN(new_n922));
  MUX2_X1   g0722(.A(new_n683), .B(new_n637), .S(new_n922), .Z(new_n923));
  OAI211_X1 g0723(.A(new_n917), .B(new_n920), .C1(new_n782), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n554), .A2(new_n668), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n567), .A2(new_n925), .A3(new_n576), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n554), .A2(new_n566), .A3(new_n668), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n671), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT44), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n671), .A2(new_n929), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT45), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n665), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n930), .B(KEYINPUT44), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT45), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n933), .B(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n666), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n657), .A2(KEYINPUT107), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n664), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n721), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n675), .B(KEYINPUT41), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n780), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n660), .A2(new_n928), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n567), .B1(new_n926), .B2(new_n493), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n669), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n948), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n923), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n666), .A2(new_n928), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n924), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT110), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(KEYINPUT110), .B(new_n924), .C1(new_n946), .C2(new_n955), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n958), .A2(new_n960), .ZN(G387));
  NOR2_X1   g0761(.A1(new_n275), .A2(G50), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT50), .ZN(new_n963));
  NAND2_X1  g0763(.A1(G68), .A2(G77), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n963), .A2(new_n296), .A3(new_n674), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n918), .B1(new_n238), .B2(new_n286), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n674), .A2(new_n728), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n213), .A2(new_n206), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n736), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n761), .A2(new_n909), .B1(new_n741), .B2(new_n905), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G311), .B2(new_n770), .ZN(new_n972));
  INV_X1    g0772(.A(G322), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n744), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  INV_X1    g0775(.A(G283), .ZN(new_n976));
  INV_X1    g0776(.A(G294), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n975), .B1(new_n976), .B2(new_n811), .C1(new_n977), .C2(new_n757), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT49), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n751), .A2(G326), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n303), .B1(new_n749), .B2(G116), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G159), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n744), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n811), .A2(new_n329), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G150), .B2(new_n751), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n246), .B2(new_n757), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n345), .B(new_n989), .C1(G97), .C2(new_n749), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G68), .A2(new_n774), .B1(new_n770), .B2(new_n395), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(new_n202), .C2(new_n741), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n984), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n734), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n781), .C1(new_n663), .C2(new_n782), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n721), .A2(new_n942), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n675), .B1(new_n721), .B2(new_n942), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n995), .B1(new_n779), .B2(new_n943), .C1(new_n997), .C2(new_n998), .ZN(G393));
  INV_X1    g0799(.A(new_n940), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n997), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n676), .B1(new_n940), .B2(new_n996), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n780), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n737), .B1(new_n214), .B2(new_n506), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n251), .B2(new_n723), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n760), .A2(new_n741), .B1(new_n744), .B2(new_n905), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT52), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n761), .A2(new_n977), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n772), .B1(new_n973), .B2(new_n750), .C1(new_n811), .C2(new_n218), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n345), .B1(new_n976), .B2(new_n757), .C1(new_n762), .C2(new_n909), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  AOI21_X1  g0813(.A(new_n345), .B1(new_n758), .B2(G68), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n388), .B2(new_n748), .C1(new_n806), .C2(new_n750), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT112), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n754), .A2(G77), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G50), .A2(new_n770), .B1(new_n774), .B2(new_n395), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n272), .A2(new_n744), .B1(new_n741), .B2(new_n985), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1006), .B1(new_n1023), .B2(new_n734), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n781), .C1(new_n782), .C2(new_n929), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1003), .A2(new_n1004), .A3(new_n1025), .ZN(G390));
  AND3_X1   g0826(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n844), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT38), .B1(new_n842), .B2(new_n844), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT39), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n845), .A2(new_n850), .A3(new_n871), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n880), .C2(new_n870), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n791), .A2(G330), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n718), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n876), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n870), .B1(new_n845), .B2(new_n850), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n689), .A2(new_n651), .A3(new_n791), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(new_n879), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1035), .B1(new_n1037), .B2(new_n876), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1031), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1032), .A2(new_n821), .A3(new_n855), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT114), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n855), .B1(new_n1032), .B2(new_n821), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1034), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1033), .A2(new_n876), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n1040), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n877), .A2(new_n879), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1045), .A2(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n366), .A2(G330), .A3(new_n453), .A4(new_n821), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n623), .C1(new_n454), .C2(new_n699), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT114), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1031), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n870), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n851), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n876), .B1(new_n1036), .B2(new_n879), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n872), .A2(new_n873), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n878), .B1(new_n698), .B2(new_n791), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1056), .B1(new_n1061), .B2(new_n876), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1054), .B(new_n1055), .C1(new_n1063), .C2(new_n1041), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1043), .A2(new_n1053), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT115), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1063), .B2(new_n1041), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n676), .B1(new_n1068), .B2(new_n1052), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1043), .A2(new_n1064), .A3(KEYINPUT115), .A4(new_n1053), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n206), .A2(new_n762), .B1(new_n761), .B2(new_n506), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n218), .A2(new_n741), .B1(new_n744), .B2(new_n976), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1017), .B1(new_n388), .B2(new_n757), .C1(new_n977), .C2(new_n750), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n345), .B1(new_n748), .B2(new_n222), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT117), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n811), .A2(new_n985), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n758), .A2(G150), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT53), .ZN(new_n1080));
  INV_X1    g0880(.A(G128), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1081), .A2(new_n744), .B1(new_n741), .B2(new_n809), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G125), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n303), .B1(new_n750), .B2(new_n1084), .C1(new_n202), .C2(new_n748), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT54), .B(G143), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n774), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1087), .C1(new_n803), .C2(new_n762), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1077), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n784), .B1(new_n1089), .B2(new_n734), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n732), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n275), .B2(new_n816), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1068), .A2(new_n780), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n780), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(G378));
  OAI21_X1  g0899(.A(new_n1052), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1051), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n859), .B(G330), .C1(new_n864), .C2(KEYINPUT40), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n883), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT56), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n279), .A2(new_n650), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n617), .A2(new_n327), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n323), .B2(new_n328), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT55), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT55), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(KEYINPUT56), .A3(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1103), .A2(new_n874), .A3(new_n875), .A4(new_n882), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1105), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1119), .B1(new_n1105), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1102), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1102), .B(KEYINPUT57), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n675), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n780), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n295), .B(new_n345), .C1(new_n757), .C2(new_n246), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n749), .A2(G58), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n976), .B2(new_n750), .C1(new_n811), .C2(new_n222), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G107), .C2(new_n742), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G97), .A2(new_n770), .B1(new_n774), .B2(new_n600), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n218), .C2(new_n744), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT58), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n202), .B1(new_n343), .B2(G41), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1137), .C1(KEYINPUT118), .C2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n770), .A2(G132), .B1(new_n758), .B2(new_n1086), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G137), .B2(new_n774), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n744), .A2(new_n1084), .B1(new_n272), .B2(new_n811), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n1081), .C2(new_n741), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G33), .B1(new_n749), .B2(G159), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n751), .B2(G124), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1139), .B(new_n1150), .C1(KEYINPUT118), .C2(new_n1138), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1151), .A2(new_n734), .B1(new_n202), .B2(new_n816), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1119), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n781), .B(new_n1152), .C1(new_n1153), .C2(new_n732), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1128), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1127), .A2(new_n1156), .ZN(G375));
  NAND2_X1  g0957(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n945), .A3(new_n1053), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1049), .A2(new_n779), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n876), .A2(new_n731), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G128), .A2(new_n751), .B1(new_n754), .B2(G50), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n985), .B2(new_n757), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n345), .B(new_n1165), .C1(G137), .C2(new_n742), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n745), .A2(G132), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT123), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G150), .A2(new_n774), .B1(new_n770), .B2(new_n1086), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1130), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n345), .B1(new_n748), .B2(new_n246), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT121), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n987), .B(new_n1172), .C1(G294), .C2(new_n745), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n909), .A2(new_n750), .B1(new_n757), .B2(new_n205), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT122), .Z(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G107), .B2(new_n774), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n742), .A2(G283), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n770), .A2(G116), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1170), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n734), .B1(new_n222), .B2(new_n816), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1163), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1162), .B1(new_n781), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1161), .A2(new_n1183), .ZN(G381));
  NOR4_X1   g0984(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(G375), .A2(G384), .A3(G378), .A4(G381), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(G407));
  INV_X1    g0987(.A(G378), .ZN(new_n1188));
  INV_X1    g0988(.A(G343), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(G213), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1156), .A3(new_n1127), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT124), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(G407), .A2(G213), .A3(new_n1194), .A4(new_n1195), .ZN(G409));
  INV_X1    g0996(.A(new_n945), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1105), .A2(new_n1120), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1153), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1105), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1200));
  AOI221_X4 g1000(.A(new_n1197), .B1(new_n1100), .B2(new_n1101), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1071), .B(new_n1098), .C1(new_n1201), .C2(new_n1155), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT125), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1128), .B(new_n1154), .C1(new_n1123), .C2(new_n1197), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1071), .A4(new_n1098), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1127), .A2(G378), .A3(new_n1156), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1053), .A2(KEYINPUT60), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n676), .B1(new_n1160), .B2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1049), .A2(KEYINPUT60), .A3(new_n1051), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT126), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT126), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1214), .A2(G384), .A3(new_n1183), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G384), .B1(new_n1214), .B2(new_n1183), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1208), .A2(new_n1190), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT62), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1208), .A2(new_n1190), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(G2897), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1214), .A2(new_n1183), .ZN(new_n1224));
  INV_X1    g1024(.A(G384), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1214), .A2(G384), .A3(new_n1183), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1221), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1220), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1208), .A2(new_n1232), .A3(new_n1190), .A4(new_n1217), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1219), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n958), .B2(new_n960), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G390), .B(new_n924), .C1(new_n946), .C2(new_n955), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(G393), .B(G396), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n956), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1237), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1238), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT127), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1245), .B(new_n1238), .C1(new_n1241), .C2(new_n1237), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1234), .A2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1247), .A2(new_n1231), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1208), .A2(KEYINPUT63), .A3(new_n1190), .A4(new_n1217), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1220), .B2(new_n1229), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1218), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1250), .B(new_n1251), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1255), .ZN(G405));
  NAND2_X1  g1056(.A1(new_n1247), .A2(new_n1217), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G375), .A2(new_n1188), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1240), .B1(new_n1216), .B2(new_n1215), .C1(new_n1244), .C2(new_n1246), .ZN(new_n1259));
  AND4_X1   g1059(.A1(new_n1207), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1257), .A2(new_n1259), .B1(new_n1258), .B2(new_n1207), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G402));
endmodule


