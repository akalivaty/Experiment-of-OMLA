//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n541, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n577, new_n580, new_n582, new_n583, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1085;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT67), .ZN(G160));
  AND2_X1   g048(.A1(new_n460), .A2(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n470), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n470), .ZN(new_n485));
  XOR2_X1   g060(.A(KEYINPUT68), .B(KEYINPUT4), .Z(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g062(.A1(KEYINPUT68), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(new_n460), .A3(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n460), .A2(new_n462), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n470), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n487), .A2(new_n491), .A3(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT69), .A2(G651), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G62), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n505), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n501), .A2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n498), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  OAI221_X1 g096(.A(new_n513), .B1(new_n514), .B2(new_n507), .C1(new_n520), .C2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n516), .ZN(new_n527));
  INV_X1    g102(.A(new_n507), .ZN(new_n528));
  AOI22_X1  g103(.A1(G52), .A2(new_n527), .B1(new_n528), .B2(G90), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT72), .B(G43), .Z(new_n533));
  OAI22_X1  g108(.A1(new_n532), .A2(new_n507), .B1(new_n516), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT73), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n527), .A2(G53), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G91), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n537), .B1(new_n507), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G299));
  NAND2_X1  g128(.A1(new_n527), .A2(G49), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n528), .A2(G87), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(G288));
  NAND3_X1  g132(.A1(new_n498), .A2(G48), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(G86), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n558), .B1(new_n507), .B2(new_n559), .C1(new_n560), .C2(new_n537), .ZN(G305));
  NAND2_X1  g136(.A1(new_n528), .A2(G85), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n527), .A2(G47), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n537), .C2(new_n564), .ZN(G290));
  NAND2_X1  g140(.A1(G301), .A2(G868), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n527), .A2(G54), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n498), .A2(G92), .A3(new_n505), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT10), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT75), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n566), .B1(new_n574), .B2(G868), .ZN(G284));
  OAI21_X1  g150(.A(new_n566), .B1(new_n574), .B2(G868), .ZN(G321));
  NAND2_X1  g151(.A1(G286), .A2(G868), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(G868), .B2(new_n552), .ZN(G297));
  OAI21_X1  g153(.A(new_n577), .B1(G868), .B2(new_n552), .ZN(G280));
  INV_X1    g154(.A(G559), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n574), .B1(new_n580), .B2(G860), .ZN(G148));
  NAND2_X1  g156(.A1(new_n574), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G868), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(G868), .B2(new_n539), .ZN(G323));
  XNOR2_X1  g159(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g160(.A1(new_n459), .A2(G2105), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n474), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n587), .B(new_n588), .Z(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT13), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(G2100), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n476), .A2(G123), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n479), .A2(G135), .ZN(new_n593));
  NOR2_X1   g168(.A1(G99), .A2(G2105), .ZN(new_n594));
  OAI21_X1  g169(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G2096), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n591), .A2(new_n598), .ZN(G156));
  XNOR2_X1  g174(.A(KEYINPUT15), .B(G2435), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT77), .B(G2438), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g177(.A(G2427), .B(G2430), .Z(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n605));
  XOR2_X1   g180(.A(G2443), .B(G2446), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(G2451), .B(G2454), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT78), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT16), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n607), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(G1341), .B(G1348), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT79), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT80), .ZN(new_n615));
  INV_X1    g190(.A(G14), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n611), .B2(new_n613), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(G401));
  XOR2_X1   g194(.A(G2084), .B(G2090), .Z(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(G2067), .B(G2678), .Z(new_n622));
  XOR2_X1   g197(.A(G2072), .B(G2078), .Z(new_n623));
  NOR3_X1   g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT81), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT18), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(KEYINPUT17), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n627), .A2(new_n622), .A3(new_n620), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT82), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n623), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n621), .B(new_n630), .C1(new_n627), .C2(new_n622), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(new_n597), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G227));
  XNOR2_X1  g210(.A(G1971), .B(G1976), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT83), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT19), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1956), .B(G2474), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT84), .ZN(new_n641));
  XOR2_X1   g216(.A(G1961), .B(G1966), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT20), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n641), .A2(new_n642), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n639), .A2(new_n643), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n645), .B(new_n648), .C1(new_n646), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G1986), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1991), .B(G1996), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT22), .B(G1981), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G229));
  INV_X1    g232(.A(G16), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G19), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n539), .B2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G1341), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(G22), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(G166), .B2(new_n658), .ZN(new_n663));
  INV_X1    g238(.A(G1971), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(G16), .A2(G23), .ZN(new_n666));
  INV_X1    g241(.A(G288), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n667), .B2(G16), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT33), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  MUX2_X1   g245(.A(G6), .B(G305), .S(G16), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT32), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n665), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT34), .ZN(new_n677));
  MUX2_X1   g252(.A(G24), .B(G290), .S(G16), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT87), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AOI22_X1  g255(.A1(G119), .A2(new_n476), .B1(new_n479), .B2(G131), .ZN(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n682));
  NOR2_X1   g257(.A1(G95), .A2(G2105), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT86), .Z(new_n684));
  OAI21_X1  g259(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(G25), .B(new_n685), .S(G29), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT35), .B(G1991), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(KEYINPUT90), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n677), .A2(new_n680), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n661), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G4), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n574), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT92), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT91), .B(G1348), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G5), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G171), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT93), .B(G2067), .Z(new_n701));
  INV_X1    g276(.A(KEYINPUT28), .ZN(new_n702));
  INV_X1    g277(.A(G26), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n476), .A2(G128), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n479), .A2(G140), .ZN(new_n707));
  NOR2_X1   g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n705), .B1(new_n710), .B2(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n704), .B1(new_n711), .B2(new_n702), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n700), .A2(G1961), .B1(new_n701), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n696), .B2(new_n697), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n693), .A2(new_n698), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT29), .B(G2090), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n586), .A2(G103), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n723), .C1(new_n470), .C2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G33), .B(new_n725), .S(G29), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2072), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n715), .A2(new_n720), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n700), .A2(G1961), .ZN(new_n730));
  NAND2_X1  g305(.A1(G160), .A2(G29), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n716), .B1(new_n732), .B2(G34), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n730), .B1(G2084), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G2084), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n716), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n716), .ZN(new_n744));
  MUX2_X1   g319(.A(new_n743), .B(new_n744), .S(KEYINPUT97), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G2078), .ZN(new_n746));
  AOI22_X1  g321(.A1(G129), .A2(new_n476), .B1(new_n479), .B2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n586), .A2(G105), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT95), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT26), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n658), .A2(KEYINPUT23), .A3(G20), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n757));
  INV_X1    g332(.A(G20), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n552), .C2(new_n658), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n755), .B(new_n761), .C1(new_n753), .C2(new_n754), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n742), .B(new_n762), .C1(new_n691), .C2(new_n692), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n745), .A2(G2078), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G21), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G168), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT96), .B(G1966), .Z(new_n768));
  XOR2_X1   g343(.A(new_n767), .B(new_n768), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n712), .A2(new_n701), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT30), .B(G28), .Z(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(G29), .B2(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n763), .A2(new_n765), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n596), .A2(new_n716), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n728), .A2(new_n729), .A3(new_n773), .A4(new_n774), .ZN(G150));
  INV_X1    g350(.A(G150), .ZN(G311));
  NAND2_X1  g351(.A1(G80), .A2(G543), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n502), .A2(new_n504), .ZN(new_n778));
  INV_X1    g353(.A(G67), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G651), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT99), .ZN(new_n782));
  AOI22_X1  g357(.A1(G55), .A2(new_n527), .B1(new_n528), .B2(G93), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G860), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT37), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n574), .A2(G559), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT39), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n784), .B(KEYINPUT100), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(new_n539), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G860), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g371(.A(KEYINPUT106), .B(G37), .ZN(new_n797));
  INV_X1    g372(.A(new_n491), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n492), .A2(new_n493), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G2105), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n485), .A2(new_n486), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n752), .B(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n710), .B(KEYINPUT102), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n725), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n685), .B(new_n589), .ZN(new_n809));
  INV_X1    g384(.A(G130), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n475), .A2(KEYINPUT104), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n479), .A2(G142), .ZN(new_n812));
  OR2_X1    g387(.A1(G106), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT104), .B1(new_n475), .B2(new_n810), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n809), .B(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n725), .A2(new_n806), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n805), .A2(new_n807), .A3(new_n818), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n808), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n808), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT105), .ZN(new_n823));
  XNOR2_X1  g398(.A(G160), .B(G162), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n596), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n797), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n822), .A2(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g407(.A(new_n790), .B(new_n582), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n552), .B(new_n573), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT41), .Z(new_n835));
  AND2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT42), .ZN(new_n839));
  XNOR2_X1  g414(.A(G303), .B(G288), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G305), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G290), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT42), .B1(new_n836), .B2(new_n838), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n839), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n839), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(G868), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n784), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g424(.A(new_n847), .B1(G868), .B2(new_n848), .ZN(G331));
  XNOR2_X1  g425(.A(G171), .B(G286), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n790), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n790), .A2(new_n851), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n837), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n835), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n842), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n790), .B(new_n851), .ZN(new_n858));
  INV_X1    g433(.A(new_n835), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n843), .A3(new_n854), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n797), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n857), .B2(new_n861), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n843), .B1(new_n860), .B2(new_n854), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n863), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT43), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n870), .B1(new_n862), .B2(new_n863), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT44), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n862), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT108), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n866), .A2(new_n880), .A3(new_n864), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n869), .B1(new_n876), .B2(new_n882), .ZN(G397));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G164), .B2(G1384), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n466), .A2(new_n471), .A3(G40), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n889), .A2(G1986), .A3(G290), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(G1986), .A3(G290), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT110), .Z(new_n893));
  XOR2_X1   g468(.A(new_n710), .B(G2067), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n752), .B(G1996), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n685), .B(new_n687), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1384), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n802), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT50), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT116), .B(G2084), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n909), .A3(new_n886), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n802), .A2(KEYINPUT45), .A3(new_n902), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n885), .A2(new_n886), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n912), .A2(KEYINPUT115), .A3(new_n768), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT115), .B1(new_n912), .B2(new_n768), .ZN(new_n914));
  OAI211_X1 g489(.A(G168), .B(new_n910), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G8), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT51), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(KEYINPUT118), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n912), .A2(new_n768), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT115), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n912), .A2(KEYINPUT115), .A3(new_n768), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n910), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(G8), .A3(G286), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n915), .B(new_n918), .C1(KEYINPUT118), .C2(new_n917), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT62), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT119), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n921), .A2(new_n928), .A3(new_n929), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n885), .B2(new_n911), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT45), .B1(new_n802), .B2(new_n902), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n886), .B1(new_n938), .B2(KEYINPUT111), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n664), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G2090), .ZN(new_n941));
  NOR3_X1   g516(.A1(G164), .A2(new_n904), .A3(G1384), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT50), .B1(new_n802), .B2(new_n902), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n941), .B(new_n886), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n916), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G303), .A2(G8), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT55), .Z(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(KEYINPUT112), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n907), .A2(new_n951), .A3(new_n941), .A4(new_n886), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n940), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n947), .A3(G8), .ZN(new_n954));
  NAND2_X1  g529(.A1(G305), .A2(G1981), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n560), .A2(new_n537), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n528), .A2(G86), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT113), .B(G1981), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n558), .A4(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(KEYINPUT49), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(KEYINPUT49), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G164), .A2(G1384), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n916), .B1(new_n965), .B2(new_n886), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n955), .A2(new_n960), .A3(new_n959), .A4(KEYINPUT49), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(G288), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n966), .B(new_n972), .C1(new_n969), .C2(G288), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n949), .A2(new_n954), .A3(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(G164), .A2(new_n884), .A3(G1384), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT111), .B1(new_n976), .B2(new_n938), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n887), .B1(new_n885), .B2(new_n936), .ZN(new_n978));
  INV_X1    g553(.A(G2078), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n907), .A2(new_n886), .ZN(new_n982));
  INV_X1    g557(.A(G1961), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n912), .A2(new_n981), .A3(G2078), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n975), .A2(G301), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n935), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT122), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n932), .B1(new_n931), .B2(new_n934), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n935), .A2(KEYINPUT122), .A3(new_n987), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n980), .A2(new_n981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n982), .A2(new_n983), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(G301), .A3(new_n996), .A4(new_n985), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT121), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT120), .B(G2078), .Z(new_n999));
  OR3_X1    g574(.A1(new_n912), .A2(new_n981), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G171), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n984), .A2(new_n1003), .A3(G301), .A4(new_n985), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT54), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n984), .A2(G301), .A3(new_n1000), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1007), .B(new_n1008), .C1(new_n986), .C2(G301), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n975), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n931), .A2(new_n934), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n552), .B(KEYINPUT57), .ZN(new_n1012));
  INV_X1    g587(.A(G1956), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n982), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n977), .A2(new_n978), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n887), .A2(new_n903), .A3(G2067), .ZN(new_n1019));
  INV_X1    g594(.A(G1348), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n982), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n573), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1017), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1021), .A2(new_n573), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT60), .B1(new_n1024), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(KEYINPUT61), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT61), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1012), .A2(new_n1027), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT60), .ZN(new_n1029));
  INV_X1    g604(.A(new_n573), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .A4(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n937), .A2(new_n939), .A3(G1996), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT58), .B(G1341), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n965), .B2(new_n886), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n539), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT59), .Z(new_n1037));
  OAI21_X1  g612(.A(new_n1023), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1010), .A2(new_n1011), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n916), .B1(new_n926), .B2(new_n910), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1040), .A2(new_n954), .A3(new_n974), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(G168), .A4(new_n949), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1040), .A2(new_n954), .A3(new_n974), .A4(G168), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n1045), .B2(new_n948), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n947), .B1(new_n953), .B2(G8), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n1045), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n974), .A2(G8), .A3(new_n947), .A4(new_n953), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n968), .A2(new_n969), .A3(new_n667), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n959), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n966), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n1039), .A2(new_n1050), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n901), .B1(new_n994), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n888), .B1(new_n895), .B2(new_n752), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT125), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n889), .A2(G1996), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT46), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  NOR2_X1   g637(.A1(new_n685), .A2(new_n687), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT123), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n897), .B2(new_n889), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(G2067), .B2(new_n710), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1066), .B(KEYINPUT124), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n888), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n890), .B(KEYINPUT126), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT48), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n900), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1062), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT127), .B1(new_n1056), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n901), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n935), .A2(KEYINPUT122), .A3(new_n987), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT122), .B1(new_n935), .B2(new_n987), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n991), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1039), .A2(new_n1050), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT127), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1072), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1073), .A2(new_n1082), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g658(.A(G401), .B(G227), .C1(new_n829), .C2(new_n830), .ZN(new_n1085));
  NAND4_X1  g659(.A1(new_n656), .A2(new_n867), .A3(G319), .A4(new_n1085), .ZN(G225));
  INV_X1    g660(.A(G225), .ZN(G308));
endmodule


