//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n219), .A2(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n220), .B2(new_n219), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n217), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n246), .A2(new_n221), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G1), .B2(new_n222), .ZN(new_n248));
  MUX2_X1   g0048(.A(new_n245), .B(new_n248), .S(G50), .Z(new_n249));
  NAND2_X1  g0049(.A1(new_n203), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n222), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n246), .A2(new_n221), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n264), .B1(new_n208), .B2(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT64), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT64), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G33), .A3(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n221), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n278), .A2(new_n270), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n279), .B2(G226), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G200), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G190), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n261), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT10), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT12), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n245), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n244), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n287), .B(G68), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G68), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n247), .B(KEYINPUT70), .C1(G1), .C2(new_n222), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(KEYINPUT12), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n291), .B(new_n294), .C1(new_n287), .C2(new_n245), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT73), .B1(new_n253), .B2(new_n202), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n255), .A2(G77), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n296), .B(new_n297), .C1(new_n222), .C2(G68), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n253), .A2(KEYINPUT73), .A3(new_n202), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n258), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT11), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT13), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n304), .A2(new_n306), .A3(G232), .A4(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(G226), .A4(new_n263), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n268), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n313), .A3(new_n268), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n272), .B1(new_n279), .B2(G238), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n310), .A2(new_n313), .A3(new_n268), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n310), .B2(new_n268), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n303), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n302), .B1(new_n322), .B2(G190), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(new_n260), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n281), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n283), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n286), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G169), .B1(new_n317), .B2(new_n321), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT14), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n327), .B1(new_n337), .B2(new_n320), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(G179), .A3(new_n320), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n302), .ZN(new_n343));
  INV_X1    g0143(.A(new_n268), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n304), .A2(new_n306), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT65), .B(G107), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT66), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n351), .B2(new_n350), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n272), .B1(new_n279), .B2(G244), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(KEYINPUT67), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT67), .B1(new_n353), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n329), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT68), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n254), .B1(new_n359), .B2(new_n253), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n359), .B2(new_n253), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT15), .B(G87), .Z(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n258), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n289), .A2(new_n290), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n208), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n293), .B2(new_n208), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n353), .A2(new_n354), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n327), .A3(new_n355), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n358), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(G190), .B1(new_n356), .B2(new_n357), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(G200), .A3(new_n355), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n371), .B1(new_n366), .B2(new_n367), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT71), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n333), .A2(new_n343), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT78), .ZN(new_n388));
  INV_X1    g0188(.A(new_n245), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n254), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n248), .B2(new_n254), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n262), .B2(G20), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n305), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT7), .B(new_n222), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n292), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  OR3_X1    g0199(.A1(new_n253), .A2(KEYINPUT74), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G58), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n292), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n201), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT74), .B1(new_n253), .B2(new_n399), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n392), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n247), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n392), .B(new_n408), .C1(new_n398), .C2(new_n405), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n391), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n304), .A2(new_n306), .A3(G226), .A4(G1698), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n304), .A2(new_n306), .A3(G223), .A4(new_n263), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n268), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n278), .A2(G232), .A3(new_n270), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT76), .ZN(new_n417));
  INV_X1    g0217(.A(new_n272), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n278), .A2(new_n419), .A3(G232), .A4(new_n270), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n415), .A2(new_n417), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n272), .B1(new_n414), .B2(new_n268), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n423), .A2(G190), .A3(new_n417), .A4(new_n420), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n388), .B(KEYINPUT17), .C1(new_n410), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n388), .A2(KEYINPUT17), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n388), .A2(KEYINPUT17), .ZN(new_n428));
  AND4_X1   g0228(.A1(new_n410), .A2(new_n427), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n409), .A3(new_n258), .ZN(new_n432));
  INV_X1    g0232(.A(new_n391), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n421), .A2(new_n327), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G179), .B2(new_n421), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT18), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n410), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT77), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(new_n437), .A3(KEYINPUT18), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n410), .B2(new_n436), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n430), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n387), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT82), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT81), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT81), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n448), .B(new_n449), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  AOI211_X1 g0255(.A(G1), .B(new_n455), .C1(new_n452), .C2(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n459));
  AOI21_X1  g0259(.A(G41), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n448), .ZN(new_n461));
  OAI211_X1 g0261(.A(G257), .B(new_n278), .C1(new_n457), .C2(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n460), .A2(new_n448), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(G274), .A3(new_n454), .A4(new_n456), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n304), .A2(new_n306), .A3(G244), .A4(new_n263), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n262), .A2(new_n468), .A3(G244), .A4(new_n263), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n304), .A2(new_n306), .A3(G250), .A4(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n344), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n467), .B2(new_n469), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT80), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n268), .B1(new_n478), .B2(KEYINPUT79), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n470), .A2(KEYINPUT79), .A3(new_n474), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n329), .B(new_n465), .C1(new_n480), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT6), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n486), .A2(new_n210), .A3(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(G97), .B(G107), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n489), .A2(new_n222), .B1(new_n208), .B2(new_n253), .ZN(new_n490));
  INV_X1    g0290(.A(new_n348), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n394), .B2(new_n397), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n258), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n389), .A2(new_n210), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n258), .B1(new_n244), .B2(G33), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n389), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n465), .B1(new_n482), .B2(new_n481), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n327), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n485), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n462), .A2(new_n464), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n477), .B2(new_n479), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(G190), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n483), .B1(new_n481), .B2(new_n482), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n477), .A2(KEYINPUT80), .A3(new_n479), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n324), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(G87), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n262), .A2(new_n222), .A3(G68), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n256), .A2(new_n210), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(KEYINPUT19), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n309), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(new_n515), .B2(KEYINPUT19), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G87), .A2(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n491), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n258), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n362), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n369), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n511), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n262), .A2(G238), .A3(new_n263), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n265), .C2(new_n209), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n268), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n455), .A2(new_n271), .A3(G1), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n529));
  INV_X1    g0329(.A(G250), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n244), .B2(G45), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(new_n529), .B1(new_n278), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n526), .A2(G190), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n327), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n497), .A2(new_n362), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n519), .A2(new_n538), .A3(new_n521), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n539), .C1(G179), .C2(new_n534), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n502), .A2(new_n510), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n502), .A2(new_n510), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT84), .ZN(new_n546));
  OAI211_X1 g0346(.A(G270), .B(new_n278), .C1(new_n457), .C2(new_n461), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n262), .A2(G257), .A3(new_n263), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n262), .A2(G264), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n347), .A2(G303), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n551), .A2(new_n552), .A3(new_n268), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n551), .B2(new_n268), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n464), .B(new_n547), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n289), .A2(G116), .A3(new_n290), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n472), .B(new_n222), .C1(G33), .C2(new_n210), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT20), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  AOI22_X1  g0359(.A1(KEYINPUT86), .A2(new_n558), .B1(new_n559), .B2(G20), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n560), .A3(new_n258), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n496), .A2(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n561), .A2(new_n562), .B1(new_n369), .B2(new_n559), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n327), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(new_n566), .A3(KEYINPUT21), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n555), .A2(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n555), .A2(new_n566), .A3(KEYINPUT87), .A4(KEYINPUT21), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n553), .A2(new_n554), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n547), .A2(new_n464), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n564), .A2(new_n565), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n574), .A2(G179), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n569), .A2(new_n572), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n265), .A2(new_n211), .B1(new_n252), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n347), .A2(new_n530), .A3(G1698), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n268), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G264), .B(new_n278), .C1(new_n457), .C2(new_n461), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n329), .A3(new_n464), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n464), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n327), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n262), .A2(new_n222), .A3(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n262), .A2(new_n590), .A3(new_n222), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n593), .A2(G107), .B1(G20), .B2(new_n524), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n491), .A2(G20), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(KEYINPUT23), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT24), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT24), .B1(new_n592), .B2(new_n596), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n597), .A2(new_n598), .A3(new_n247), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n495), .A2(G107), .A3(new_n245), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT88), .ZN(new_n601));
  INV_X1    g0401(.A(G107), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n244), .A2(new_n602), .A3(G13), .A4(G20), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n603), .A2(new_n601), .A3(new_n604), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT89), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n585), .B(new_n587), .C1(new_n599), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n598), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n592), .A2(new_n596), .A3(KEYINPUT24), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n258), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n586), .A2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT89), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n609), .B(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n582), .A2(new_n583), .A3(new_n464), .A4(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n614), .A2(new_n615), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n576), .B1(new_n555), .B2(G200), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n574), .A2(G190), .A3(new_n575), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n578), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n447), .A2(new_n544), .A3(new_n546), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n611), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n619), .B1(new_n578), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n545), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n502), .B2(new_n541), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n542), .A2(new_n501), .A3(new_n485), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n540), .B(KEYINPUT90), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n447), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n438), .A2(new_n440), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n358), .A2(new_n377), .A3(new_n373), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n325), .B1(new_n342), .B2(new_n302), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n426), .A2(new_n429), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n331), .B1(new_n640), .B2(new_n286), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(G369));
  AND2_X1   g0442(.A1(new_n222), .A2(G13), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n244), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(G343), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n576), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n578), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n578), .A2(new_n623), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n650), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n611), .A2(new_n649), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n649), .B1(new_n599), .B2(new_n610), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n619), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n611), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n655), .ZN(new_n664));
  INV_X1    g0464(.A(new_n649), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n578), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n663), .A2(new_n664), .A3(new_n668), .ZN(G399));
  NAND3_X1  g0469(.A1(new_n491), .A2(new_n559), .A3(new_n517), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n218), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n224), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n665), .B1(new_n628), .B2(new_n633), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(KEYINPUT29), .B(new_n665), .C1(new_n628), .C2(new_n633), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n555), .A2(new_n329), .ZN(new_n683));
  INV_X1    g0483(.A(new_n534), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n584), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n685), .A3(new_n505), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n683), .A2(new_n685), .A3(KEYINPUT30), .A4(new_n505), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n555), .A2(new_n329), .A3(new_n534), .A4(new_n586), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n688), .B(new_n689), .C1(new_n509), .C2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n649), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n546), .A2(new_n624), .A3(new_n544), .A4(new_n665), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n691), .B2(new_n649), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n682), .A2(new_n697), .A3(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT92), .B1(new_n682), .B2(new_n697), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n677), .B1(new_n702), .B2(G1), .ZN(G364));
  AOI21_X1  g0503(.A(new_n244), .B1(new_n643), .B2(G45), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n673), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n654), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G330), .B2(new_n653), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n262), .A2(new_n218), .ZN(new_n709));
  INV_X1    g0509(.A(G355), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n710), .B1(G116), .B2(new_n218), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n239), .A2(new_n455), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n672), .A2(new_n262), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n455), .B2(new_n225), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n711), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n221), .B1(G20), .B2(new_n327), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n706), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n329), .A2(new_n324), .ZN(new_n724));
  AND2_X1   g0524(.A1(G20), .A2(G190), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G326), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n324), .A2(G179), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n725), .ZN(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n726), .A2(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n329), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n725), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n262), .B(new_n731), .C1(G322), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n222), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT33), .B(G317), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n728), .A2(new_n736), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(G283), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n736), .A2(new_n732), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G329), .A2(new_n745), .B1(new_n746), .B2(G311), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n222), .B1(new_n743), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G294), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n735), .A2(new_n742), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n726), .A2(new_n202), .B1(new_n733), .B2(new_n401), .ZN(new_n752));
  INV_X1    g0552(.A(new_n746), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n753), .A2(new_n208), .B1(new_n292), .B2(new_n737), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n752), .B(new_n754), .C1(G97), .C2(new_n749), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n744), .A2(new_n399), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT93), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT32), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(KEYINPUT32), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G87), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n262), .B1(new_n729), .B2(new_n761), .C1(new_n602), .C2(new_n740), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n751), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n765));
  INV_X1    g0565(.A(new_n720), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n764), .B2(KEYINPUT95), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n723), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n719), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n653), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n708), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  NAND2_X1  g0572(.A1(new_n373), .A2(new_n649), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n382), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n378), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n637), .A2(new_n665), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n678), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n378), .A2(new_n649), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n774), .B2(new_n378), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n780), .B(new_n665), .C1(new_n628), .C2(new_n633), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n706), .B1(new_n782), .B2(new_n697), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n697), .B2(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(new_n706), .ZN(new_n785));
  INV_X1    g0585(.A(G137), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n726), .A2(new_n786), .B1(new_n737), .B2(new_n251), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT98), .ZN(new_n788));
  INV_X1    g0588(.A(G143), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n789), .B2(new_n733), .C1(new_n399), .C2(new_n753), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT34), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n262), .B1(new_n740), .B2(new_n292), .ZN(new_n792));
  INV_X1    g0592(.A(G132), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n729), .A2(new_n202), .B1(new_n744), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(G58), .C2(new_n749), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n738), .A2(G283), .B1(new_n746), .B2(G116), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n740), .A2(new_n761), .B1(new_n744), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT97), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n347), .B1(new_n726), .B2(new_n730), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n602), .A2(new_n729), .B1(new_n733), .B2(new_n579), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G97), .C2(new_n749), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n798), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n766), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n720), .A2(new_n717), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n785), .B(new_n806), .C1(new_n208), .C2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT99), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n718), .B2(new_n780), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n784), .A2(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n489), .ZN(new_n812));
  OAI211_X1 g0612(.A(G116), .B(new_n223), .C1(new_n812), .C2(KEYINPUT35), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(KEYINPUT35), .B2(new_n812), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n225), .B(G77), .C1(new_n401), .C2(new_n292), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n202), .A2(G68), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n244), .B(G13), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n341), .B1(new_n338), .B2(new_n339), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n334), .A2(KEYINPUT14), .ZN(new_n821));
  OAI211_X1 g0621(.A(KEYINPUT100), .B(new_n302), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT100), .B1(new_n342), .B2(new_n302), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n823), .A2(new_n824), .A3(new_n649), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n410), .A2(new_n647), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n446), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT101), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n446), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n434), .A2(new_n437), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n410), .A2(new_n425), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n834), .B2(new_n827), .ZN(new_n835));
  INV_X1    g0635(.A(new_n827), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n832), .A4(new_n833), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n829), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n839), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n828), .B2(KEYINPUT101), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n831), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n826), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n827), .B1(new_n639), .B2(new_n635), .ZN(new_n847));
  OAI211_X1 g0647(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n834), .C2(new_n827), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(KEYINPUT102), .C2(new_n839), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n841), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n845), .A2(new_n850), .A3(new_n826), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n825), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n636), .A2(new_n648), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n781), .A2(new_n776), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n302), .A2(new_n649), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n325), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n823), .B2(new_n824), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n342), .A2(new_n302), .A3(new_n649), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n842), .A2(new_n845), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT103), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n447), .A2(new_n680), .A3(new_n681), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n641), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n865), .B(new_n867), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n845), .A2(new_n850), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n777), .B1(new_n857), .B2(new_n858), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n870), .A2(new_n696), .A3(KEYINPUT40), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n696), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n842), .B2(new_n845), .ZN(new_n874));
  OAI211_X1 g0674(.A(G330), .B(new_n872), .C1(new_n874), .C2(KEYINPUT40), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n447), .A2(G330), .A3(new_n696), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n870), .A2(new_n696), .ZN(new_n877));
  AND4_X1   g0677(.A1(KEYINPUT38), .A2(new_n829), .A3(new_n831), .A4(new_n839), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n844), .B2(new_n831), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(new_n881), .B1(new_n869), .B2(new_n871), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n447), .A2(new_n696), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n875), .A2(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n868), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n244), .B2(new_n643), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n868), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n819), .B1(new_n886), .B2(new_n887), .ZN(G367));
  INV_X1    g0688(.A(KEYINPUT111), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n668), .A2(new_n664), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n502), .A2(new_n665), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n502), .A2(new_n510), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n503), .A2(new_n649), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT45), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT44), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n663), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n663), .B1(new_n896), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n653), .A2(G330), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n666), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(new_n658), .Z(new_n905));
  AOI21_X1  g0705(.A(new_n701), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n673), .B(KEYINPUT41), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n704), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n892), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT105), .B1(new_n668), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT105), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n658), .A2(new_n667), .A3(new_n912), .A4(new_n892), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n510), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n502), .B1(new_n917), .B2(new_n611), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n665), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(KEYINPUT42), .A3(new_n913), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n665), .A2(new_n522), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n632), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n542), .A2(new_n922), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n916), .A2(new_n926), .A3(new_n919), .A4(new_n920), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n663), .A2(new_n894), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n937), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n939), .A2(new_n934), .B1(new_n663), .B2(new_n894), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n909), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G97), .A2(new_n741), .B1(new_n746), .B2(G283), .ZN(new_n942));
  INV_X1    g0742(.A(G317), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n744), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n726), .A2(new_n799), .B1(new_n733), .B2(new_n730), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT107), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n347), .B1(new_n737), .B2(new_n579), .C1(new_n491), .C2(new_n748), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n729), .A2(new_n559), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  OR4_X1    g0749(.A1(new_n944), .A2(new_n946), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n738), .A2(G159), .B1(new_n746), .B2(G50), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n729), .A2(new_n401), .B1(new_n744), .B2(new_n786), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT109), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n262), .B1(new_n733), .B2(new_n251), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n726), .A2(new_n789), .B1(new_n740), .B2(new_n208), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(G68), .C2(new_n749), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n952), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT110), .Z(new_n960));
  AOI21_X1  g0760(.A(new_n766), .B1(new_n960), .B2(KEYINPUT47), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT47), .B2(new_n960), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n235), .A2(new_n714), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n722), .B1(new_n672), .B2(new_n362), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n785), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n962), .B(new_n965), .C1(new_n769), .C2(new_n930), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n889), .B1(new_n941), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n940), .A2(new_n938), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n896), .A2(new_n899), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n661), .A3(new_n662), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n663), .A2(new_n896), .A3(new_n899), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n904), .B(new_n658), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n702), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n705), .B1(new_n974), .B2(new_n907), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n889), .B(new_n966), .C1(new_n968), .C2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(G387));
  OAI21_X1  g0779(.A(new_n905), .B1(new_n699), .B2(new_n700), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n682), .A2(new_n697), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT92), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n698), .A3(new_n973), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n984), .A3(new_n673), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n658), .A2(new_n769), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n713), .B1(new_n232), .B2(new_n455), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n671), .B2(new_n709), .ZN(new_n988));
  AOI21_X1  g0788(.A(G45), .B1(G68), .B2(G77), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n254), .A2(KEYINPUT50), .A3(G50), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT50), .B1(new_n254), .B2(G50), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n671), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n988), .A2(new_n992), .B1(new_n602), .B2(new_n672), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n706), .B1(new_n993), .B2(new_n722), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n729), .A2(new_n208), .B1(new_n744), .B2(new_n251), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n347), .B(new_n995), .C1(G97), .C2(new_n741), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n753), .A2(new_n292), .B1(new_n399), .B2(new_n726), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n737), .A2(new_n254), .B1(new_n733), .B2(new_n202), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n996), .B(new_n999), .C1(new_n520), .C2(new_n748), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n726), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n1001), .A2(G322), .B1(new_n746), .B2(G303), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n799), .B2(new_n737), .C1(new_n943), .C2(new_n733), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT112), .Z(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n729), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G294), .A2(new_n1007), .B1(new_n749), .B2(G283), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n262), .B1(new_n745), .B2(G326), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n559), .C2(new_n740), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1000), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n994), .B1(new_n1015), .B2(new_n720), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n905), .A2(new_n705), .B1(new_n986), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n985), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT113), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n985), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(G393));
  INV_X1    g0822(.A(new_n980), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n902), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n972), .A2(new_n980), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n1025), .A3(new_n673), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n894), .A2(new_n719), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n737), .A2(new_n730), .B1(new_n748), .B2(new_n559), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT114), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(G294), .B2(new_n746), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT115), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G283), .A2(new_n1007), .B1(new_n745), .B2(G322), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n347), .C1(new_n602), .C2(new_n740), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT52), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n726), .A2(new_n943), .B1(new_n733), .B2(new_n799), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1032), .B(new_n1037), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n737), .A2(new_n202), .B1(new_n729), .B2(new_n292), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n726), .A2(new_n251), .B1(new_n733), .B2(new_n399), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT51), .Z(new_n1041));
  OAI22_X1  g0841(.A1(new_n753), .A2(new_n254), .B1(new_n744), .B2(new_n789), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n262), .B1(new_n748), .B2(new_n208), .C1(new_n761), .C2(new_n740), .ZN(new_n1043));
  OR4_X1    g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n766), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n242), .A2(new_n714), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n722), .B(new_n1046), .C1(G97), .C2(new_n672), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n785), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n902), .A2(new_n705), .B1(new_n1027), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1026), .A2(new_n1049), .ZN(G390));
  INV_X1    g0850(.A(new_n859), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n697), .B2(new_n777), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n870), .A2(new_n696), .A3(G330), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n854), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n866), .A2(new_n876), .A3(new_n641), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n854), .A3(new_n1053), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n825), .B1(new_n854), .B2(new_n859), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n845), .A2(new_n850), .A3(new_n826), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n825), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n860), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n869), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1053), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1066), .B1(new_n846), .B2(new_n851), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1061), .A2(new_n845), .A3(new_n850), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1053), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1060), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1068), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n1071), .A3(new_n1053), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n1059), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n673), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n785), .B1(new_n254), .B2(new_n807), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1001), .A2(G283), .B1(new_n746), .B2(G97), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n491), .B2(new_n737), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT117), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n733), .A2(new_n559), .B1(new_n748), .B2(new_n208), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT118), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n347), .B1(new_n729), .B2(new_n761), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n740), .A2(new_n292), .B1(new_n744), .B2(new_n579), .ZN(new_n1087));
  NOR4_X1   g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT54), .B(G143), .Z(new_n1089));
  AOI22_X1  g0889(.A1(new_n738), .A2(G137), .B1(new_n746), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT116), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G128), .A2(new_n1001), .B1(new_n741), .B2(G50), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n744), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n729), .A2(new_n251), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT53), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n262), .C1(new_n793), .C2(new_n733), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1095), .A2(new_n1096), .B1(new_n399), .B2(new_n748), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1094), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1081), .A2(new_n1088), .B1(new_n1091), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1078), .B1(new_n1101), .B2(new_n766), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n846), .A2(new_n851), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n717), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n705), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1077), .A2(new_n1106), .ZN(G378));
  AOI21_X1  g0907(.A(new_n1065), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n853), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n878), .A2(new_n879), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n860), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n882), .B(G330), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n286), .A2(new_n332), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT55), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n260), .A2(new_n648), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n875), .A2(new_n852), .A3(new_n863), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1118), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n705), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(G33), .A2(G41), .ZN(new_n1123));
  AOI211_X1 g0923(.A(G50), .B(new_n1123), .C1(new_n347), .C2(new_n449), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n449), .B(new_n347), .C1(new_n729), .C2(new_n208), .ZN(new_n1125));
  INV_X1    g0925(.A(G283), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n740), .A2(new_n401), .B1(new_n744), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G68), .C2(new_n749), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G116), .A2(new_n1001), .B1(new_n734), .B2(G107), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n738), .A2(G97), .B1(new_n746), .B2(new_n362), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT58), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n737), .A2(new_n793), .B1(new_n733), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1007), .A2(new_n1089), .B1(new_n746), .B2(G137), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1093), .B2(new_n726), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G150), .C2(new_n749), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT59), .Z(new_n1139));
  OR2_X1    g0939(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n745), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n1123), .C1(new_n399), .C2(new_n740), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1133), .B1(new_n1132), .B2(new_n1131), .C1(new_n1139), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n720), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n785), .B1(new_n202), .B2(new_n807), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1118), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1146), .C1(new_n1147), .C2(new_n718), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1122), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n866), .A2(new_n876), .A3(new_n641), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1059), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1120), .A2(new_n1121), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n673), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1147), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1112), .A2(new_n1119), .A3(new_n1118), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1073), .A2(new_n1057), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1149), .B1(new_n1154), .B2(new_n1160), .ZN(G375));
  AND3_X1   g0961(.A1(new_n1052), .A2(new_n854), .A3(new_n1053), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n854), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1150), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n1059), .A3(new_n907), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n785), .B1(new_n292), .B2(new_n807), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n729), .A2(new_n399), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n753), .A2(new_n251), .B1(new_n744), .B2(new_n1134), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n738), .C2(new_n1089), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n262), .B1(new_n740), .B2(new_n401), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n726), .A2(new_n793), .B1(new_n733), .B2(new_n786), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G50), .C2(new_n749), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n753), .A2(new_n491), .B1(new_n579), .B2(new_n726), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n737), .A2(new_n559), .B1(new_n744), .B2(new_n730), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n347), .B1(new_n740), .B2(new_n208), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n210), .A2(new_n729), .B1(new_n733), .B2(new_n1126), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n362), .C2(new_n749), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1169), .A2(new_n1172), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1166), .B1(new_n1179), .B2(new_n766), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1051), .B2(new_n717), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n705), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1165), .A2(new_n1183), .ZN(G381));
  NOR2_X1   g0984(.A1(G390), .A2(G381), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n978), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1159), .B(KEYINPUT57), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n673), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G378), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1149), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1019), .A2(new_n771), .A3(new_n1021), .ZN(new_n1193));
  OR3_X1    g0993(.A1(new_n1193), .A2(KEYINPUT121), .A3(G384), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT121), .B1(new_n1193), .B2(G384), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1186), .A2(KEYINPUT122), .A3(new_n1192), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n978), .A2(new_n1196), .A3(new_n1185), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1191), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(G407));
  AND2_X1   g1001(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1202));
  INV_X1    g1002(.A(G213), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1191), .A2(new_n1203), .A3(G343), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT123), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1203), .A2(G343), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1192), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT124), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT124), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(G407), .A2(new_n1212), .A3(new_n1209), .A4(new_n1206), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(G409));
  NAND2_X1  g1014(.A1(new_n1207), .A2(G2897), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1057), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n673), .B(new_n1059), .C1(new_n1216), .C2(KEYINPUT60), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1164), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G384), .B(new_n1183), .C1(new_n1217), .C2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1216), .A2(KEYINPUT60), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1164), .A2(new_n1218), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n673), .A4(new_n1059), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G384), .B1(new_n1224), .B2(new_n1183), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1215), .B1(new_n1221), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1183), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1227));
  INV_X1    g1027(.A(G384), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1215), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1220), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1226), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1221), .A2(new_n1225), .A3(new_n1215), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1229), .B2(new_n1220), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT125), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1190), .B1(new_n1189), .B2(new_n1149), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1122), .A2(new_n1077), .A3(new_n1106), .A4(new_n1148), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1152), .A2(new_n908), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1238), .A2(new_n1239), .B1(new_n1203), .B2(G343), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1233), .B(new_n1236), .C1(new_n1237), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT63), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G375), .A2(G378), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1239), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1207), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n941), .A2(new_n966), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n985), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1020), .B1(new_n985), .B2(new_n1017), .ZN(new_n1254));
  OAI21_X1  g1054(.A(G396), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1193), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n1256), .B2(KEYINPUT111), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1255), .A2(new_n1193), .B1(new_n1026), .B2(new_n1049), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1252), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(G390), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n889), .B1(new_n1255), .B2(new_n1193), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1251), .C1(G390), .C2(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1250), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT126), .B1(new_n1249), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1240), .B1(G378), .B2(G375), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1241), .A2(KEYINPUT63), .B1(new_n1244), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1265), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1260), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1248), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1248), .B2(new_n1275), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1274), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1267), .A2(new_n1271), .B1(new_n1272), .B2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(new_n1243), .A2(new_n1191), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1244), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1272), .ZN(G402));
endmodule


