//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(new_n205), .B2(new_n206), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT23), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  INV_X1    g019(.A(new_n214), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT67), .B(G176gat), .Z(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(G169gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT23), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n219), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n209), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n208), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n230), .A2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n208), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n223), .B1(new_n236), .B2(KEYINPUT25), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(KEYINPUT1), .B2(new_n238), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT27), .B(G183gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT28), .A3(new_n206), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT70), .Z(new_n252));
  NOR3_X1   g051(.A1(new_n205), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n205), .A2(KEYINPUT69), .ZN(new_n254));
  AOI211_X1 g053(.A(G190gat), .B(new_n253), .C1(KEYINPUT27), .C2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(KEYINPUT28), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n214), .A2(new_n257), .A3(new_n215), .ZN(new_n258));
  OAI221_X1 g057(.A(new_n258), .B1(new_n257), .B2(new_n214), .C1(new_n205), .C2(new_n206), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n237), .A2(new_n249), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n249), .B1(new_n237), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n203), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n266));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n237), .A2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n248), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n202), .B1(new_n271), .B2(new_n262), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(KEYINPUT33), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n202), .A3(new_n262), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT34), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT34), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n271), .A2(new_n276), .A3(new_n202), .A4(new_n262), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n277), .ZN(new_n279));
  INV_X1    g078(.A(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n265), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n266), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT31), .B(G50gat), .ZN(new_n285));
  INV_X1    g084(.A(G106gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G141gat), .B(G148gat), .Z(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT2), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(new_n294), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  AND2_X1   g099(.A1(G211gat), .A2(G218gat), .ZN(new_n301));
  AND2_X1   g100(.A1(G197gat), .A2(G204gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G197gat), .A2(G204gat), .ZN(new_n303));
  OAI22_X1  g102(.A1(KEYINPUT22), .A2(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n305), .B2(new_n304), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n309), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n300), .A3(new_n297), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G228gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n308), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n310), .B2(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT82), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n300), .B1(new_n323), .B2(KEYINPUT82), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n298), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT83), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n329), .B(new_n298), .C1(new_n325), .C2(new_n326), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n322), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(G22gat), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n323), .A2(KEYINPUT82), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(new_n300), .A3(new_n324), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n329), .B1(new_n334), .B2(new_n298), .ZN(new_n335));
  INV_X1    g134(.A(new_n330), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n321), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G22gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n318), .B(KEYINPUT81), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G78gat), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n332), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n288), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n332), .A2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G78gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n287), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n279), .A2(new_n282), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n350));
  INV_X1    g149(.A(new_n266), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n284), .A2(new_n344), .A3(new_n348), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n312), .ZN(new_n354));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n355), .B(KEYINPUT74), .Z(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n270), .B2(new_n314), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n237), .B2(new_n261), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n270), .A2(new_n356), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n237), .B2(new_n261), .ZN(new_n361));
  INV_X1    g160(.A(new_n355), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n312), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  NAND4_X1  g165(.A1(new_n359), .A2(KEYINPUT30), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n359), .B2(new_n363), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT75), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(new_n363), .A3(new_n366), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n359), .A2(KEYINPUT76), .A3(new_n363), .A4(new_n366), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XOR2_X1   g177(.A(G57gat), .B(G85gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n299), .A2(new_n249), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n298), .A2(new_n248), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n298), .A2(new_n248), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n248), .A3(new_n313), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n394), .A2(new_n381), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n393), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n382), .B2(new_n399), .ZN(new_n404));
  INV_X1    g203(.A(new_n381), .ZN(new_n405));
  INV_X1    g204(.A(new_n396), .ZN(new_n406));
  NOR4_X1   g205(.A1(new_n404), .A2(KEYINPUT5), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n380), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n380), .A3(new_n408), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n359), .A2(new_n363), .ZN(new_n416));
  INV_X1    g215(.A(new_n366), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n367), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n370), .A2(new_n376), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT35), .B1(new_n353), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n344), .A2(new_n348), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n351), .B1(new_n349), .B2(new_n350), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n368), .A2(new_n369), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n376), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n380), .B(KEYINPUT85), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n386), .A2(new_n389), .B1(new_n397), .B2(new_n400), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n407), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n433), .A3(new_n410), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT35), .B1(new_n434), .B2(new_n412), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n423), .A2(new_n426), .A3(new_n429), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n422), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n382), .A2(new_n381), .A3(new_n383), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(KEYINPUT86), .A3(KEYINPUT39), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n430), .C1(KEYINPUT39), .C2(new_n438), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n448), .A2(new_n433), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n416), .B2(KEYINPUT37), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n359), .A2(KEYINPUT87), .A3(new_n363), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n357), .A2(new_n358), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(new_n312), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n360), .B(new_n354), .C1(new_n362), .C2(new_n361), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n417), .A3(new_n459), .ZN(new_n460));
  AND4_X1   g259(.A1(new_n412), .A2(new_n373), .A3(new_n434), .A4(new_n375), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n366), .B1(new_n452), .B2(new_n454), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n416), .A2(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n450), .B(new_n423), .C1(new_n462), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n424), .B2(new_n425), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n284), .A2(KEYINPUT36), .A3(new_n352), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n344), .A2(new_n348), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n469), .A2(new_n470), .B1(new_n421), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n472), .B2(KEYINPUT84), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n421), .A2(new_n471), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n437), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G15gat), .B(G22gat), .Z(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G1gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(G1gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT16), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n483));
  INV_X1    g282(.A(G8gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n484), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n489));
  INV_X1    g288(.A(G29gat), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT14), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n494), .C1(G29gat), .C2(G36gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G43gat), .B(G50gat), .Z(new_n498));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT88), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n493), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT14), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n497), .A2(new_n500), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT14), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n508));
  OAI211_X1 g307(.A(KEYINPUT15), .B(new_n501), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT17), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  AOI211_X1 g314(.A(new_n483), .B(new_n484), .C1(new_n479), .C2(new_n482), .ZN(new_n516));
  INV_X1    g315(.A(new_n487), .ZN(new_n517));
  AND4_X1   g316(.A1(new_n517), .A2(new_n479), .A3(new_n482), .A4(new_n485), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n509), .B(new_n506), .C1(new_n516), .C2(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(KEYINPUT91), .A3(new_n524), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n519), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n515), .B(KEYINPUT13), .Z(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n515), .A4(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G197gat), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT11), .B(G169gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT12), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT92), .B1(new_n530), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n523), .A2(new_n528), .A3(new_n535), .A4(new_n529), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n477), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(new_n290), .ZN(new_n547));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(G57gat), .A2(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(G57gat), .A2(G64gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G127gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n557), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n558), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n519), .B1(KEYINPUT21), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n565), .A2(new_n566), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n567), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n567), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n550), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n575), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n578), .A3(new_n549), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(KEYINPUT7), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n596), .A2(new_n592), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n590), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n599), .B2(new_n602), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n604), .A2(new_n513), .A3(new_n512), .A4(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n603), .A2(new_n510), .B1(KEYINPUT41), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n607), .B2(new_n610), .ZN(new_n614));
  OR3_X1    g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n612), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT96), .Z(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n615), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(KEYINPUT101), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n585), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G120gat), .B(G148gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT104), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT105), .Z(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G230gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n317), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n561), .B1(new_n599), .B2(new_n602), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n601), .A2(new_n600), .A3(new_n590), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n597), .A2(new_n598), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n574), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(KEYINPUT102), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n603), .A2(new_n640), .A3(new_n574), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(new_n644), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n639), .B2(new_n641), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n643), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n634), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n642), .A2(new_n634), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n631), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n631), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT106), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n651), .A2(new_n657), .A3(new_n653), .A4(new_n631), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n626), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n545), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n415), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n481), .ZN(G1324gat));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n545), .A2(new_n428), .A3(new_n661), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(G8gat), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT42), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n665), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n672), .A2(KEYINPUT107), .A3(new_n674), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(new_n662), .ZN(new_n679));
  AOI21_X1  g478(.A(G15gat), .B1(new_n679), .B2(new_n426), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT108), .ZN(new_n681));
  INV_X1    g480(.A(new_n474), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n679), .B2(new_n683), .ZN(G1326gat));
  AND2_X1   g483(.A1(new_n545), .A2(new_n471), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n661), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n622), .A2(new_n624), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n639), .A2(new_n641), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT103), .B1(new_n691), .B2(KEYINPUT10), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n646), .B1(new_n649), .B2(new_n643), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n652), .B1(new_n694), .B2(new_n634), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n657), .B1(new_n695), .B2(new_n631), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n633), .B1(new_n692), .B2(new_n693), .ZN(new_n697));
  INV_X1    g496(.A(new_n631), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n652), .A4(new_n698), .ZN(new_n699));
  OAI22_X1  g498(.A1(new_n696), .A2(new_n699), .B1(new_n695), .B2(new_n631), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n690), .A2(new_n700), .A3(new_n585), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n545), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n415), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n490), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n477), .A2(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n472), .A2(new_n467), .B1(new_n422), .B2(new_n436), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n709), .B2(new_n690), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n541), .B(KEYINPUT93), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT109), .B1(new_n539), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n543), .B(new_n714), .C1(new_n538), .C2(new_n537), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n700), .A2(new_n585), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n711), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n415), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n720), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n491), .A3(new_n428), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n719), .B2(new_n429), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(G43gat), .B1(new_n719), .B2(new_n474), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n702), .A2(new_n727), .A3(new_n426), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT110), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n719), .B2(new_n423), .ZN(new_n732));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n685), .A2(new_n733), .A3(new_n701), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n735), .B(new_n736), .Z(G1331gat));
  NOR4_X1   g536(.A1(new_n709), .A2(new_n625), .A3(new_n659), .A4(new_n717), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n703), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n428), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n682), .ZN(new_n745));
  INV_X1    g544(.A(new_n426), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(G71gat), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n745), .A2(G71gat), .B1(new_n738), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n471), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n467), .A2(new_n472), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n690), .B1(new_n752), .B2(new_n437), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n717), .A2(new_n585), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT113), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(KEYINPUT51), .A3(new_n754), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n703), .A2(new_n700), .A3(new_n594), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT114), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n717), .A2(new_n585), .A3(new_n659), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n711), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(new_n703), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n594), .B2(new_n765), .ZN(G1336gat));
  NOR3_X1   g565(.A1(new_n429), .A2(G92gat), .A3(new_n659), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n756), .B2(new_n758), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n708), .A2(new_n428), .A3(new_n710), .A4(new_n763), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(new_n769), .B2(G92gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n757), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n767), .B1(new_n773), .B2(new_n755), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n775), .B2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n777), .B(new_n778), .C1(new_n772), .C2(new_n774), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n771), .B(KEYINPUT116), .C1(new_n776), .C2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1337gat));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n682), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G99gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n759), .A2(new_n700), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n746), .A2(G99gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(G1338gat));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n764), .A2(new_n471), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT117), .B(G106gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n423), .A2(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n790), .B(new_n793), .C1(new_n787), .C2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n700), .B(new_n794), .C1(new_n773), .C2(new_n755), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n790), .B2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n625), .B1(new_n713), .B2(new_n715), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n659), .ZN(new_n802));
  AND4_X1   g601(.A1(new_n800), .A2(new_n716), .A3(new_n626), .A4(new_n659), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n631), .B1(new_n697), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n692), .A2(new_n693), .A3(new_n633), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n656), .A2(new_n658), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n808), .A3(KEYINPUT55), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n527), .B1(new_n525), .B2(new_n526), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n515), .B1(new_n514), .B2(new_n520), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n534), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n543), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n814), .A2(new_n690), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n659), .B2(new_n818), .ZN(new_n821));
  INV_X1    g620(.A(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n700), .A2(new_n822), .A3(KEYINPUT119), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n821), .B(new_n823), .C1(new_n716), .C2(new_n814), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n824), .B2(new_n690), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n804), .B1(new_n825), .B2(new_n585), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n703), .ZN(new_n827));
  INV_X1    g626(.A(new_n353), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n429), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT120), .Z(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n717), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n428), .A2(new_n415), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n826), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n544), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(G1340gat));
  NAND3_X1  g636(.A1(new_n830), .A2(new_n243), .A3(new_n700), .ZN(new_n838));
  OAI21_X1  g637(.A(G120gat), .B1(new_n834), .B2(new_n659), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1341gat));
  INV_X1    g639(.A(new_n585), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n834), .A2(new_n566), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n566), .B1(new_n829), .B2(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n843), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1342gat));
  OR3_X1    g646(.A1(new_n829), .A2(G134gat), .A3(new_n690), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n834), .B2(new_n690), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  AND2_X1   g651(.A1(new_n474), .A2(new_n833), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n826), .B2(new_n471), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n471), .A2(KEYINPUT57), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n544), .A2(new_n812), .A3(new_n811), .A4(new_n813), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n700), .A2(new_n822), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n689), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n841), .B1(new_n858), .B2(new_n819), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n804), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n853), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G141gat), .B1(new_n861), .B2(new_n835), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n682), .A2(new_n423), .A3(new_n428), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n835), .A2(G141gat), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT124), .Z(new_n867));
  OAI211_X1 g666(.A(new_n862), .B(new_n863), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT122), .B(new_n853), .C1(new_n854), .C2(new_n860), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n717), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n872), .B2(G141gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n865), .A2(new_n867), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n868), .B1(new_n876), .B2(new_n863), .ZN(G1344gat));
  OAI21_X1  g676(.A(new_n859), .B1(new_n544), .B2(new_n660), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(new_n471), .ZN(new_n879));
  INV_X1    g678(.A(new_n826), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n879), .A2(KEYINPUT57), .B1(new_n880), .B2(new_n855), .ZN(new_n881));
  XOR2_X1   g680(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n882));
  NOR2_X1   g681(.A1(new_n659), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n853), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n870), .A2(new_n871), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n659), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(KEYINPUT59), .ZN(new_n887));
  INV_X1    g686(.A(new_n865), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n700), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n882), .A2(G148gat), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n887), .A2(G148gat), .B1(new_n889), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n885), .B2(new_n841), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(new_n290), .A3(new_n585), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  NOR3_X1   g693(.A1(new_n885), .A2(new_n291), .A3(new_n690), .ZN(new_n895));
  AOI21_X1  g694(.A(G162gat), .B1(new_n888), .B2(new_n689), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n429), .A2(new_n703), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n353), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n826), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n835), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n717), .A2(new_n225), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(G1348gat));
  INV_X1    g703(.A(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n700), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(new_n224), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT126), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(KEYINPUT126), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n908), .B(new_n909), .C1(new_n213), .C2(new_n906), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n585), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n205), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n250), .B2(new_n911), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT60), .Z(G1350gat));
  OAI22_X1  g713(.A1(new_n901), .A2(new_n690), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n682), .A2(new_n899), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n881), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n835), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n826), .A2(new_n471), .A3(new_n918), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n717), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n920), .B2(new_n926), .ZN(G1352gat));
  OAI21_X1  g726(.A(G204gat), .B1(new_n919), .B2(new_n659), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n922), .A2(G204gat), .A3(new_n659), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  NOR2_X1   g730(.A1(new_n841), .A2(G211gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n924), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n881), .A2(new_n585), .A3(new_n918), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n919), .B2(new_n690), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n690), .A2(G218gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n925), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1355gat));
endmodule


