//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053;
  AND2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G155gat), .B(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT2), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G113gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT68), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G113gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(G120gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G134gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G127gat), .ZN(new_n230));
  INV_X1    g029(.A(G127gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G134gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(G120gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n232), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(KEYINPUT3), .A2(new_n220), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n220), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n234), .B1(new_n227), .B2(new_n225), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n238), .A2(new_n233), .B1(new_n230), .B2(new_n232), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n220), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n242), .A2(new_n245), .B1(new_n248), .B2(KEYINPUT4), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n251), .A3(new_n241), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n252), .A3(new_n243), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT84), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(KEYINPUT84), .A3(new_n258), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT39), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n236), .A2(new_n241), .B1(new_n219), .B2(new_n209), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(new_n257), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267));
  AOI211_X1 g066(.A(new_n267), .B(new_n257), .C1(new_n249), .C2(new_n255), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G1gat), .B(G29gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT40), .A4(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n258), .B1(new_n248), .B2(new_n263), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n236), .A2(new_n241), .A3(new_n219), .A4(new_n209), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n220), .B1(new_n246), .B2(new_n247), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n257), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n253), .A2(new_n286), .A3(KEYINPUT4), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n253), .B2(KEYINPUT4), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n279), .A2(KEYINPUT4), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n258), .B1(new_n242), .B2(new_n245), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n249), .A2(new_n255), .A3(new_n282), .A4(new_n257), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n274), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n269), .A3(new_n274), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT40), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G211gat), .A2(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n299), .B(new_n306), .C1(new_n303), .C2(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G226gat), .ZN(new_n311));
  INV_X1    g110(.A(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT23), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(KEYINPUT23), .B2(new_n317), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT24), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT66), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(KEYINPUT65), .A3(new_n332), .ZN(new_n333));
  OR3_X1    g132(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n327), .A2(new_n331), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n332), .ZN(new_n337));
  NAND3_X1  g136(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n330), .ZN(new_n339));
  INV_X1    g138(.A(G169gat), .ZN(new_n340));
  INV_X1    g139(.A(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT64), .B1(new_n342), .B2(new_n319), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n317), .A2(new_n316), .A3(KEYINPUT23), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n339), .B(new_n323), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n324), .A2(new_n335), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n342), .B1(new_n322), .B2(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n317), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n325), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G183gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n354), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n329), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n352), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n362), .A2(new_n352), .A3(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n351), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n315), .B1(new_n346), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n336), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n335), .A2(KEYINPUT25), .A3(new_n321), .A4(new_n323), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(KEYINPUT67), .ZN(new_n370));
  AOI21_X1  g169(.A(G190gat), .B1(new_n357), .B2(new_n354), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT28), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n325), .B(new_n350), .C1(new_n372), .C2(new_n363), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n373), .A3(KEYINPUT74), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n314), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n346), .B2(new_n365), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n310), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n366), .A2(new_n376), .A3(new_n374), .ZN(new_n380));
  INV_X1    g179(.A(new_n310), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n369), .A2(new_n373), .A3(new_n313), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n379), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n388), .A2(KEYINPUT76), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT76), .B1(new_n388), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n383), .A4(new_n387), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n386), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT75), .B(new_n387), .C1(new_n379), .C2(new_n383), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n275), .B(new_n298), .C1(new_n392), .C2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n310), .B1(new_n245), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G228gat), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(new_n312), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n310), .A2(new_n404), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n243), .B1(new_n408), .B2(new_n244), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n308), .B2(new_n309), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n410), .B(new_n220), .C1(new_n412), .C2(KEYINPUT3), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n407), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n309), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n300), .A2(new_n302), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT73), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(KEYINPUT80), .A3(new_n299), .A4(new_n306), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n422), .A3(new_n308), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n404), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT81), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n426), .A3(new_n404), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n244), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n405), .B1(new_n428), .B2(new_n220), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n406), .A2(new_n312), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n403), .B(new_n415), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n402), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n244), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n423), .B2(new_n404), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n220), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n405), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n430), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n409), .A2(new_n410), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n413), .ZN(new_n441));
  OAI21_X1  g240(.A(G22gat), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n431), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n442), .B(new_n431), .C1(new_n432), .C2(new_n402), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n379), .A2(new_n448), .A3(new_n383), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n386), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n379), .B2(new_n383), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n447), .B(KEYINPUT38), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n346), .A2(new_n365), .A3(new_n315), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT74), .B1(new_n369), .B2(new_n373), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n313), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n381), .B1(new_n456), .B2(new_n377), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT37), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n386), .A3(new_n449), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n447), .B1(new_n460), .B2(KEYINPUT38), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n274), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n253), .A2(KEYINPUT4), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT77), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n253), .A2(new_n286), .A3(KEYINPUT4), .ZN(new_n466));
  INV_X1    g265(.A(new_n289), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n284), .B1(new_n468), .B2(new_n291), .ZN(new_n469));
  INV_X1    g268(.A(new_n294), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n288), .A2(new_n289), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n292), .B1(new_n473), .B2(new_n466), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n294), .B(new_n274), .C1(new_n474), .C2(new_n284), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT6), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n381), .B1(new_n375), .B2(new_n378), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n380), .A2(new_n310), .A3(new_n382), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(KEYINPUT37), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n449), .A3(new_n481), .A4(new_n386), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(new_n388), .A3(new_n477), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n399), .B(new_n446), .C1(new_n462), .C2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n250), .B(new_n252), .C1(new_n346), .C2(new_n365), .ZN(new_n485));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n250), .A2(new_n252), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n369), .A3(new_n373), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT32), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT33), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G15gat), .B(G43gat), .Z(new_n494));
  XNOR2_X1  g293(.A(G71gat), .B(G99gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n490), .B(KEYINPUT32), .C1(new_n492), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n489), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n486), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n487), .B1(new_n485), .B2(new_n489), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n497), .A2(new_n499), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT72), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n500), .A2(new_n509), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT71), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n500), .A2(new_n509), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n500), .B2(new_n509), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT72), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n515), .B1(new_n500), .B2(new_n509), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT36), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n476), .A2(new_n477), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n388), .A2(new_n389), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n388), .A2(KEYINPUT76), .A3(new_n389), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n393), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n386), .B1(new_n457), .B2(new_n458), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n395), .A2(new_n394), .A3(new_n386), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n446), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n519), .A2(new_n527), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n446), .A2(new_n523), .A3(new_n526), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT35), .B1(new_n542), .B2(new_n539), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n528), .A2(new_n533), .A3(new_n538), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n510), .B1(new_n524), .B2(new_n525), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n446), .A4(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n484), .A2(new_n541), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NOR3_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(KEYINPUT89), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n552));
  NOR4_X1   g351(.A1(new_n552), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G50gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT15), .B1(new_n555), .B2(G43gat), .ZN(new_n556));
  INV_X1    g355(.A(G43gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(G50gat), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  INV_X1    g358(.A(G36gat), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT88), .B(G50gat), .Z(new_n563));
  AOI21_X1  g362(.A(KEYINPUT87), .B1(new_n555), .B2(G43gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n563), .A2(new_n557), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n554), .B(new_n562), .C1(new_n567), .C2(KEYINPUT15), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n556), .A2(new_n558), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n549), .A2(KEYINPUT86), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n549), .A2(KEYINPUT86), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n550), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n559), .A2(new_n560), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n574), .A3(KEYINPUT17), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n576), .A2(G1gat), .ZN(new_n577));
  INV_X1    g376(.A(G8gat), .ZN(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT16), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT91), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n577), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT88), .B(G50gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n566), .ZN(new_n586));
  OAI22_X1  g385(.A1(G43gat), .A2(new_n585), .B1(new_n586), .B2(new_n564), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT15), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n561), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT86), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n549), .B(new_n590), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n591), .A2(new_n550), .B1(new_n559), .B2(new_n560), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n589), .A2(new_n554), .B1(new_n592), .B2(new_n569), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n575), .B(new_n584), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n584), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n568), .A2(new_n574), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n595), .A2(new_n598), .A3(KEYINPUT18), .A4(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(KEYINPUT13), .Z(new_n601));
  NOR2_X1   g400(.A1(new_n596), .A2(new_n597), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n593), .A2(new_n584), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(KEYINPUT92), .A3(new_n607), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n340), .ZN(new_n615));
  INV_X1    g414(.A(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT12), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT93), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n605), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n606), .A2(KEYINPUT92), .A3(new_n607), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT92), .B1(new_n606), .B2(new_n607), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n628));
  INV_X1    g427(.A(new_n622), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n624), .A3(new_n608), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT94), .B1(new_n548), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n519), .A2(new_n527), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n540), .A2(new_n539), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n484), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n543), .A2(new_n547), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n632), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n594), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n597), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT7), .ZN(new_n646));
  NAND2_X1  g445(.A1(G99gat), .A2(G106gat), .ZN(new_n647));
  INV_X1    g446(.A(G85gat), .ZN(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(KEYINPUT8), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G99gat), .B(G106gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n646), .B2(new_n650), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n644), .A2(new_n575), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  AND2_X1   g457(.A1(G232gat), .A2(G233gat), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G190gat), .B(G218gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n657), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n668));
  XNOR2_X1  g467(.A(G134gat), .B(G162gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n663), .B(new_n665), .C1(KEYINPUT99), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G57gat), .B(G64gat), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(G71gat), .A2(G78gat), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n676), .A2(new_n677), .B1(KEYINPUT95), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G71gat), .B(G78gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI221_X1 g481(.A(new_n680), .B1(KEYINPUT95), .B2(new_n678), .C1(new_n676), .C2(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n654), .B1(new_n651), .B2(new_n685), .ZN(new_n686));
  AOI211_X1 g485(.A(KEYINPUT100), .B(new_n652), .C1(new_n646), .C2(new_n650), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n682), .B(new_n683), .C1(new_n653), .C2(new_n655), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n682), .A2(new_n683), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT10), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n656), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(G230gat), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n690), .A2(new_n693), .B1(new_n694), .B2(new_n312), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n312), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n688), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(G120gat), .B(G148gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT101), .ZN(new_n700));
  XOR2_X1   g499(.A(G176gat), .B(G204gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n695), .A2(new_n697), .A3(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n596), .B1(KEYINPUT21), .B2(new_n684), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT96), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT21), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT96), .B1(new_n684), .B2(KEYINPUT21), .ZN(new_n714));
  AND4_X1   g513(.A1(G231gat), .A2(new_n713), .A3(G233gat), .A4(new_n714), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n713), .A2(new_n714), .B1(G231gat), .B2(G233gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  INV_X1    g517(.A(G231gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n312), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n713), .A2(G231gat), .A3(new_n714), .A4(G233gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n709), .ZN(new_n722));
  XNOR2_X1  g521(.A(G127gat), .B(G155gat), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT20), .Z(new_n724));
  AND3_X1   g523(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n717), .B2(new_n722), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n708), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n715), .A2(new_n716), .A3(new_n710), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n709), .B1(new_n720), .B2(new_n721), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n708), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n722), .A3(new_n724), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(G183gat), .B(G211gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n727), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n727), .B2(new_n734), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n675), .B(new_n707), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT102), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(KEYINPUT102), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n642), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n528), .A2(KEYINPUT103), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n528), .A2(KEYINPUT103), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g547(.A1(new_n538), .A2(new_n533), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT16), .B(G8gat), .Z(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(KEYINPUT42), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n749), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G8gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n751), .B2(new_n755), .ZN(G1325gat));
  INV_X1    g555(.A(new_n742), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n757), .A2(G15gat), .A3(new_n517), .ZN(new_n758));
  OAI21_X1  g557(.A(G15gat), .B1(new_n757), .B2(new_n635), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1326gat));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n540), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT43), .B(G22gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1327gat));
  INV_X1    g562(.A(new_n736), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n725), .A2(new_n726), .A3(new_n708), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n727), .A2(new_n734), .A3(new_n736), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n674), .A3(new_n707), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n634), .B2(new_n641), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n559), .A3(new_n746), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n671), .A2(new_n779), .A3(new_n673), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n671), .B2(new_n673), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n548), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n639), .A2(KEYINPUT44), .A3(new_n674), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT104), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n767), .A2(new_n788), .A3(new_n768), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(new_n633), .A3(new_n706), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n777), .B1(new_n793), .B2(new_n745), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G29gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n793), .A2(new_n777), .A3(new_n745), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n775), .B(new_n776), .C1(new_n795), .C2(new_n796), .ZN(G1328gat));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n560), .A3(new_n749), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n786), .A2(new_n749), .A3(new_n792), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n799), .A2(new_n800), .B1(G36gat), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n799), .A2(KEYINPUT107), .A3(new_n800), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(G1329gat));
  AND2_X1   g605(.A1(KEYINPUT108), .A2(G43gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n793), .B2(new_n635), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n772), .A2(KEYINPUT108), .A3(new_n557), .A4(new_n546), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1330gat));
  AOI21_X1  g612(.A(new_n563), .B1(new_n772), .B2(new_n540), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n446), .A2(new_n585), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n786), .A2(new_n792), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(KEYINPUT48), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT48), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(G1331gat));
  NAND4_X1  g619(.A1(new_n769), .A2(new_n633), .A3(new_n675), .A4(new_n706), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT109), .Z(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n639), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n746), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G57gat), .ZN(G1332gat));
  INV_X1    g624(.A(new_n749), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n828), .B(new_n829), .Z(G1333gat));
  INV_X1    g629(.A(G71gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n823), .A2(new_n831), .A3(new_n546), .ZN(new_n832));
  INV_X1    g631(.A(new_n635), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n834), .B2(new_n831), .ZN(new_n835));
  XOR2_X1   g634(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(G1334gat));
  NAND2_X1  g636(.A1(new_n823), .A2(new_n540), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g638(.A1(new_n769), .A2(new_n632), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n707), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n786), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G85gat), .B1(new_n843), .B2(new_n745), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n548), .B2(new_n675), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n484), .A2(new_n635), .A3(new_n636), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n546), .A2(new_n446), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n528), .A2(new_n538), .A3(new_n533), .A4(new_n545), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n523), .A2(new_n526), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n544), .A3(new_n446), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n852), .B2(KEYINPUT35), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT111), .B(new_n674), .C1(new_n847), .C2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n846), .A2(new_n840), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n846), .A2(new_n854), .A3(KEYINPUT51), .A4(new_n840), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n746), .A2(new_n648), .A3(new_n706), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n844), .B1(new_n862), .B2(new_n863), .ZN(G1336gat));
  NAND4_X1  g663(.A1(new_n784), .A2(new_n785), .A3(new_n749), .A4(new_n842), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n865), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT113), .B1(new_n865), .B2(G92gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n826), .A2(G92gat), .A3(new_n707), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n857), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n859), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n865), .B2(G92gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1337gat));
  OAI21_X1  g676(.A(G99gat), .B1(new_n843), .B2(new_n635), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n517), .A2(G99gat), .A3(new_n707), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n862), .B2(new_n879), .ZN(G1338gat));
  OR3_X1    g679(.A1(new_n446), .A2(G106gat), .A3(new_n707), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n871), .B2(new_n859), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n784), .A2(new_n785), .A3(new_n540), .A4(new_n842), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(G106gat), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n858), .A2(new_n859), .ZN(new_n886));
  INV_X1    g685(.A(new_n861), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n889));
  OR2_X1    g688(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n888), .B2(new_n890), .ZN(G1339gat));
  NOR2_X1   g690(.A1(new_n739), .A2(new_n632), .ZN(new_n892));
  INV_X1    g691(.A(new_n705), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n688), .A2(new_n689), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n692), .ZN(new_n895));
  INV_X1    g694(.A(new_n693), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n696), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n702), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n896), .A3(new_n696), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n695), .A3(KEYINPUT54), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT55), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT55), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n893), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n602), .A2(new_n603), .A3(new_n601), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n599), .B1(new_n595), .B2(new_n598), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n618), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n631), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n782), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n631), .A2(new_n706), .A3(new_n909), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n632), .B2(new_n906), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(new_n782), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n892), .B1(new_n914), .B2(new_n790), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n745), .A2(new_n749), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n848), .A3(new_n633), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n915), .A2(new_n917), .ZN(new_n920));
  INV_X1    g719(.A(new_n542), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n632), .A2(new_n222), .A3(new_n224), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n919), .A2(new_n221), .B1(new_n922), .B2(new_n923), .ZN(G1340gat));
  INV_X1    g723(.A(new_n922), .ZN(new_n925));
  AOI21_X1  g724(.A(G120gat), .B1(new_n925), .B2(new_n706), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n918), .A2(new_n848), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n707), .A2(new_n226), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G1341gat));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n231), .A3(new_n769), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n918), .A2(new_n848), .A3(new_n790), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n231), .ZN(G1342gat));
  NOR2_X1   g731(.A1(new_n918), .A2(new_n675), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n229), .A3(new_n921), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n229), .B1(new_n927), .B2(new_n674), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n935), .A2(new_n936), .ZN(G1343gat));
  NOR2_X1   g736(.A1(new_n833), .A2(new_n446), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n632), .A2(new_n210), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT116), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT117), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT117), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT58), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n916), .A2(new_n635), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n915), .B2(new_n446), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n446), .A2(new_n946), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT115), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n900), .A2(new_n695), .A3(KEYINPUT54), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n703), .B1(new_n695), .B2(KEYINPUT54), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT55), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n902), .A2(new_n949), .A3(new_n904), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n705), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n630), .A2(new_n631), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n623), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n675), .B1(new_n957), .B2(new_n912), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n769), .B1(new_n958), .B2(new_n911), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n948), .B1(new_n959), .B2(new_n892), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n945), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n210), .B1(new_n961), .B2(new_n632), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n944), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n960), .ZN(new_n965));
  INV_X1    g764(.A(new_n945), .ZN(new_n966));
  AND4_X1   g765(.A1(new_n964), .A2(new_n965), .A3(new_n632), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n964), .B1(new_n961), .B2(new_n632), .ZN(new_n968));
  OAI21_X1  g767(.A(G141gat), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n941), .B(KEYINPUT118), .Z(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT58), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(G1344gat));
  AND2_X1   g772(.A1(new_n920), .A2(new_n938), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n211), .A3(new_n706), .ZN(new_n975));
  XOR2_X1   g774(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n976));
  AND3_X1   g775(.A1(new_n741), .A2(new_n633), .A3(new_n740), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n906), .A2(new_n674), .A3(new_n910), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n769), .B1(new_n958), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n946), .B(new_n540), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT57), .B1(new_n915), .B2(new_n446), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n706), .A3(new_n966), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n976), .B1(new_n983), .B2(G148gat), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT59), .B(new_n211), .C1(new_n961), .C2(new_n706), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n975), .B1(new_n984), .B2(new_n985), .ZN(G1345gat));
  AND2_X1   g785(.A1(new_n974), .A2(new_n769), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(G155gat), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n790), .A2(new_n206), .ZN(new_n991));
  AOI22_X1  g790(.A1(new_n989), .A2(new_n990), .B1(new_n961), .B2(new_n991), .ZN(G1346gat));
  NAND3_X1  g791(.A1(new_n933), .A2(new_n207), .A3(new_n938), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT122), .ZN(new_n994));
  INV_X1    g793(.A(new_n961), .ZN(new_n995));
  OAI21_X1  g794(.A(G162gat), .B1(new_n995), .B2(new_n783), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1347gat));
  NOR4_X1   g796(.A1(new_n915), .A2(new_n826), .A3(new_n542), .A4(new_n746), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n998), .A2(new_n340), .A3(new_n632), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n745), .A2(new_n749), .A3(new_n546), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n446), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n1002), .A2(new_n1003), .A3(new_n915), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n340), .B1(new_n1004), .B2(new_n632), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n999), .B1(new_n1007), .B2(new_n1008), .ZN(G1348gat));
  NAND3_X1  g808(.A1(new_n998), .A2(new_n341), .A3(new_n706), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n1004), .A2(new_n706), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n1011), .B2(new_n341), .ZN(G1349gat));
  NAND3_X1  g811(.A1(new_n998), .A2(new_n353), .A3(new_n769), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1004), .A2(new_n791), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n1014), .B2(new_n328), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n329), .A3(new_n782), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n329), .B1(new_n1004), .B2(new_n674), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(G1351gat));
  NOR2_X1   g821(.A1(new_n915), .A2(new_n746), .ZN(new_n1023));
  NOR3_X1   g822(.A1(new_n833), .A2(new_n826), .A3(new_n446), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g824(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g825(.A(G197gat), .B1(new_n1026), .B2(new_n632), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n833), .A2(new_n746), .A3(new_n826), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n982), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n633), .A2(new_n616), .ZN(new_n1030));
  AOI21_X1  g829(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G1352gat));
  XNOR2_X1  g830(.A(KEYINPUT125), .B(G204gat), .ZN(new_n1032));
  NOR3_X1   g831(.A1(new_n1025), .A2(new_n707), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g832(.A(new_n1033), .B(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n982), .A2(new_n706), .A3(new_n1028), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1035), .A2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1034), .A2(new_n1036), .ZN(G1353gat));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1038));
  NAND4_X1  g837(.A1(new_n980), .A2(new_n769), .A3(new_n981), .A4(new_n1028), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1039), .A2(G211gat), .ZN(new_n1040));
  INV_X1    g839(.A(KEYINPUT63), .ZN(new_n1041));
  OAI21_X1  g840(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g841(.A1(new_n1039), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OR3_X1    g844(.A1(new_n1025), .A2(G211gat), .A3(new_n770), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1045), .A2(new_n1046), .ZN(G1354gat));
  INV_X1    g846(.A(G218gat), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1048), .B1(new_n1025), .B2(new_n783), .ZN(new_n1049));
  INV_X1    g848(.A(KEYINPUT127), .ZN(new_n1050));
  NOR2_X1   g849(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AND2_X1   g850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g851(.A1(new_n675), .A2(new_n1048), .ZN(new_n1053));
  AOI211_X1 g852(.A(new_n1051), .B(new_n1052), .C1(new_n1029), .C2(new_n1053), .ZN(G1355gat));
endmodule


