//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066;
  OR2_X1    g000(.A1(KEYINPUT65), .A2(G137), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT65), .A2(G137), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT11), .A2(G134), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT11), .A2(G134), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT11), .A2(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G104), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G101), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n199), .A3(G104), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n199), .A2(G104), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT79), .A2(G101), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT79), .A2(G101), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n205), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n208), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT79), .A2(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT79), .A2(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n202), .A3(new_n217), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT80), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n204), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n224), .A3(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G143), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n231), .B2(G146), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(G146), .B1(new_n222), .B2(new_n224), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(G128), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n220), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n204), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n209), .A2(new_n213), .A3(new_n205), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT80), .B1(new_n215), .B2(new_n218), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(G128), .B1(new_n226), .B2(new_n235), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n234), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n198), .B1(new_n238), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT12), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n190), .A2(new_n196), .A3(new_n193), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n196), .B1(new_n190), .B2(new_n193), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n248), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n220), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n223), .A2(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n244), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n228), .B1(new_n259), .B2(KEYINPUT1), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n247), .B1(new_n260), .B2(new_n232), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n242), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n254), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT12), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n240), .A2(new_n241), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n206), .A2(new_n208), .A3(new_n202), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G101), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n234), .B2(new_n245), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n267), .A3(G101), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n225), .A2(new_n227), .A3(new_n271), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n246), .B2(new_n247), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n270), .A2(new_n277), .B1(new_n242), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n220), .B2(new_n237), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n254), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n283), .B(new_n285), .Z(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n251), .A2(new_n265), .A3(new_n282), .A4(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n280), .A2(new_n254), .A3(new_n281), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT82), .B(G469), .Z(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n282), .B1(new_n264), .B2(new_n263), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n250), .A2(KEYINPUT12), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT81), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n251), .A2(new_n265), .A3(new_n299), .A4(new_n282), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n286), .A3(new_n300), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n289), .A2(new_n290), .A3(new_n286), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  OAI21_X1  g121(.A(G221), .B1(new_n307), .B2(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n266), .A2(new_n320), .A3(new_n204), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n318), .A2(G119), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n316), .A2(G116), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT66), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G113), .B1(new_n317), .B2(KEYINPUT5), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT66), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT66), .B1(new_n317), .B2(new_n319), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT5), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n330), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n321), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n268), .A2(G101), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n314), .A3(new_n328), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n338), .A2(new_n267), .B1(new_n339), .B2(new_n320), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n270), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n313), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n329), .A2(new_n322), .A3(new_n330), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT83), .B1(new_n334), .B2(new_n335), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n341), .B(new_n312), .C1(new_n346), .C2(new_n321), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n246), .A2(new_n349), .A3(new_n247), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n274), .B2(new_n276), .ZN(new_n351));
  INV_X1    g165(.A(G224), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G953), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n271), .A2(new_n272), .ZN(new_n356));
  INV_X1    g170(.A(new_n245), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n259), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n225), .A2(new_n227), .A3(new_n271), .ZN(new_n359));
  OAI21_X1  g173(.A(G125), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n246), .A2(new_n349), .A3(new_n247), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(new_n313), .C1(new_n337), .C2(new_n342), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n348), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n354), .A2(new_n362), .B1(KEYINPUT7), .B2(new_n353), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n353), .A2(KEYINPUT7), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n350), .B2(new_n351), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n347), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n312), .B(KEYINPUT8), .Z(new_n372));
  OAI21_X1  g186(.A(new_n320), .B1(new_n344), .B2(new_n345), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n220), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n325), .A2(new_n326), .A3(new_n323), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n242), .B(new_n320), .C1(new_n330), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n367), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n311), .B1(new_n366), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n368), .A2(new_n347), .A3(new_n370), .ZN(new_n381));
  INV_X1    g195(.A(new_n377), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n348), .A2(new_n363), .A3(new_n365), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n310), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G214), .B1(G237), .B2(G902), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n383), .A2(new_n384), .A3(new_n310), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT84), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n309), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(KEYINPUT68), .A2(G237), .ZN(new_n392));
  NOR2_X1   g206(.A1(KEYINPUT68), .A2(G237), .ZN(new_n393));
  OAI211_X1 g207(.A(G214), .B(new_n284), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n222), .A2(new_n224), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT68), .B(G237), .ZN(new_n398));
  AOI21_X1  g212(.A(G143), .B1(new_n223), .B2(new_n395), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(G214), .A3(new_n284), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G125), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(G125), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(new_n244), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT74), .B(G140), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT75), .B1(new_n409), .B2(new_n349), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT74), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G140), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n411), .B(G125), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n406), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n408), .B1(new_n416), .B2(G146), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n412), .A2(G140), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n349), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n405), .B1(new_n421), .B2(new_n411), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n244), .B1(new_n422), .B2(new_n410), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(new_n408), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n403), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n401), .A2(new_n196), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n397), .A2(G131), .A3(new_n400), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT16), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n422), .B2(new_n410), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT16), .B1(new_n404), .B2(G125), .ZN(new_n433));
  OAI21_X1  g247(.A(G146), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n435));
  INV_X1    g249(.A(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n244), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n429), .A2(new_n428), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n430), .A2(new_n434), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G113), .B(G122), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n201), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n426), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n426), .B2(new_n439), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n367), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G475), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n436), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n447), .A2(G146), .B1(new_n429), .B2(new_n427), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n416), .A2(KEYINPUT19), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT87), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n416), .A2(new_n451), .A3(KEYINPUT19), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n406), .A2(new_n407), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n450), .A2(new_n244), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n441), .B1(new_n456), .B2(new_n426), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n446), .B1(new_n457), .B2(new_n442), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n426), .A2(new_n439), .A3(new_n441), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n424), .B1(new_n423), .B2(new_n408), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n455), .A2(new_n448), .B1(new_n463), .B2(new_n403), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n460), .B1(new_n464), .B2(new_n441), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n458), .A2(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n465), .A2(KEYINPUT88), .A3(new_n459), .A4(new_n466), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n445), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(G234), .A2(G237), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(G952), .A3(new_n284), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n471), .A2(G902), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT21), .B(G898), .Z(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT93), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n318), .A2(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT14), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n318), .A3(G122), .ZN(new_n483));
  INV_X1    g297(.A(G122), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G116), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G107), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT91), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n480), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n485), .B2(new_n480), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n199), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n231), .A2(G128), .ZN(new_n494));
  INV_X1    g308(.A(G134), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n228), .A2(G143), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n494), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G134), .B1(new_n494), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n492), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(G107), .A3(new_n490), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n506), .A2(new_n493), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n488), .A2(new_n500), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT71), .B(G217), .Z(new_n509));
  NOR3_X1   g323(.A1(new_n509), .A2(G953), .A3(new_n307), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  OAI221_X1 g326(.A(new_n510), .B1(new_n504), .B2(new_n507), .C1(new_n488), .C2(new_n500), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT92), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n508), .A2(new_n515), .A3(new_n511), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n367), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n519), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n367), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n470), .A2(new_n479), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n391), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n509), .B1(G234), .B2(new_n367), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G221), .ZN(new_n528));
  INV_X1    g342(.A(G234), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n528), .A2(new_n529), .A3(G953), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT22), .B(G137), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT78), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n530), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n530), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n228), .A2(G119), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n228), .A2(G119), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n228), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G110), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n316), .A2(G128), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n550), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n550), .B2(new_n544), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G110), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n549), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR4_X1   g371(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT73), .A4(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n437), .B2(new_n434), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n244), .B1(new_n435), .B2(new_n436), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n544), .A2(new_n543), .ZN(new_n562));
  INV_X1    g376(.A(G110), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n562), .A2(new_n546), .A3(new_n563), .A4(new_n550), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n563), .A4(new_n546), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n566), .B(new_n567), .C1(new_n554), .C2(new_n556), .ZN(new_n568));
  INV_X1    g382(.A(new_n408), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n541), .B1(new_n560), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n553), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n550), .A2(new_n544), .A3(new_n551), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n556), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n554), .A2(new_n549), .A3(new_n556), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n576), .A2(new_n577), .B1(G110), .B2(new_n547), .ZN(new_n578));
  AOI211_X1 g392(.A(G146), .B(new_n433), .C1(new_n416), .C2(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n561), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n434), .A2(new_n568), .A3(new_n569), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n533), .A2(new_n530), .A3(new_n537), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n538), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n572), .A2(new_n367), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n572), .A2(new_n584), .A3(KEYINPUT25), .A4(new_n367), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n527), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n572), .A2(new_n584), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n526), .A2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n187), .A2(new_n495), .A3(new_n188), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n196), .B1(G134), .B2(G137), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n197), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n246), .B2(new_n247), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n274), .A2(new_n276), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT67), .B1(new_n254), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n357), .B1(new_n231), .B2(G146), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n603), .A2(new_n273), .B1(new_n232), .B2(new_n271), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT67), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n198), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n600), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n339), .A2(new_n320), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n608), .B(new_n600), .C1(new_n602), .C2(new_n606), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT28), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT28), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n198), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n248), .A2(new_n197), .A3(new_n598), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(new_n608), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n398), .A2(G210), .A3(new_n284), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT27), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT26), .B(G101), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n617), .A2(KEYINPUT29), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT30), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n614), .A2(new_n615), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n607), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n608), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n602), .A2(new_n606), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n609), .A3(new_n615), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n621), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT29), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n613), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n617), .A2(new_n621), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n623), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT70), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(KEYINPUT70), .A3(G472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n620), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n619), .B(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n617), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n644), .B1(new_n634), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n607), .B2(new_n609), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n648));
  INV_X1    g462(.A(new_n625), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n628), .A2(new_n615), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(KEYINPUT30), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n647), .B(new_n648), .C1(new_n651), .C2(new_n609), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n629), .A2(new_n621), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n608), .B2(new_n626), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT31), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n646), .B(new_n652), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(G472), .A2(G902), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n656), .A2(KEYINPUT32), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT32), .B1(new_n656), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n595), .B1(new_n642), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n525), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n211), .A2(new_n212), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G3));
  NAND2_X1  g479(.A1(new_n656), .A2(new_n367), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(KEYINPUT94), .A3(G472), .ZN(new_n667));
  NAND2_X1  g481(.A1(KEYINPUT94), .A2(G472), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n656), .A2(new_n367), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n594), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n309), .ZN(new_n671));
  INV_X1    g485(.A(new_n387), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n379), .B2(new_n385), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n478), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT33), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n514), .A2(new_n675), .A3(new_n516), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT33), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(G478), .A3(new_n367), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n517), .A2(new_n518), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n470), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT34), .B(G104), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G6));
  NAND3_X1  g499(.A1(new_n465), .A2(new_n459), .A3(new_n466), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n523), .B(new_n445), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n671), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT35), .B(G107), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NAND2_X1  g507(.A1(new_n667), .A2(new_n669), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n587), .A2(new_n588), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n526), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT95), .B1(new_n560), .B2(new_n571), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT95), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n580), .A2(new_n698), .A3(new_n581), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n697), .A2(new_n701), .A3(new_n699), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n591), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n696), .A2(KEYINPUT96), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT96), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n592), .B1(new_n703), .B2(new_n704), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n708), .B1(new_n589), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n694), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n391), .A2(new_n712), .A3(new_n524), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT37), .B(G110), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G12));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT96), .B1(new_n696), .B2(new_n706), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n589), .A2(new_n709), .A3(new_n708), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n308), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n251), .A2(new_n282), .A3(new_n265), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n287), .B1(new_n721), .B2(KEYINPUT81), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n302), .B1(new_n722), .B2(new_n300), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n720), .B1(new_n724), .B2(new_n295), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT97), .B(G900), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n475), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n473), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n689), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n719), .A2(new_n725), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n656), .A2(new_n657), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT32), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n656), .A2(KEYINPUT32), .A3(new_n657), .ZN(new_n738));
  INV_X1    g552(.A(G472), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n632), .B1(new_n607), .B2(new_n609), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n617), .B(new_n621), .C1(new_n740), .C2(new_n613), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n611), .B1(new_n626), .B2(new_n608), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n741), .B(new_n631), .C1(new_n742), .C2(new_n621), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n639), .B(new_n739), .C1(new_n743), .C2(new_n623), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT70), .B1(new_n637), .B2(G472), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n737), .B(new_n738), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n673), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n716), .B1(new_n734), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n379), .A2(new_n385), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n387), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n642), .B2(new_n660), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n309), .A2(new_n711), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT99), .A4(new_n733), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G128), .ZN(G30));
  NAND2_X1  g569(.A1(new_n386), .A2(new_n389), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT38), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n644), .B1(new_n627), .B2(new_n629), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n610), .A2(new_n611), .A3(new_n621), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT100), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OR3_X1    g574(.A1(new_n610), .A2(new_n611), .A3(new_n621), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT100), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n761), .B(new_n762), .C1(new_n644), .C2(new_n742), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n367), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(G472), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n737), .A3(new_n738), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n458), .A2(new_n459), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n465), .A2(new_n466), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n468), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n770), .A2(new_n445), .B1(new_n520), .B2(new_n522), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n589), .A2(new_n709), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n387), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n757), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n731), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n725), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT103), .Z(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT40), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT40), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n776), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n396), .ZN(G45));
  NAND4_X1  g599(.A1(new_n746), .A2(new_n719), .A3(new_n725), .A4(new_n673), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n470), .A2(new_n680), .A3(new_n731), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n244), .ZN(G48));
  NAND2_X1  g603(.A1(new_n288), .A2(new_n291), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n367), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT104), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n292), .A2(KEYINPUT104), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n308), .B(new_n295), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n661), .A2(new_n682), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT41), .B(G113), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G15));
  NAND4_X1  g613(.A1(new_n690), .A2(new_n796), .A3(new_n746), .A4(new_n594), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G116), .ZN(G18));
  NOR2_X1   g615(.A1(new_n795), .A2(new_n750), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n746), .A3(new_n524), .A4(new_n719), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G119), .ZN(G21));
  OAI21_X1  g618(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n621), .B1(new_n612), .B2(new_n617), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n657), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n739), .B1(new_n656), .B2(new_n367), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n595), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n673), .A2(new_n470), .A3(new_n523), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n478), .A4(new_n796), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G122), .ZN(G24));
  AND3_X1   g627(.A1(new_n470), .A2(new_n680), .A3(new_n731), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n808), .A2(new_n809), .A3(new_n773), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n802), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G125), .ZN(G27));
  INV_X1    g631(.A(KEYINPUT42), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n722), .A2(KEYINPUT105), .A3(new_n300), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT105), .B1(new_n722), .B2(new_n300), .ZN(new_n820));
  OAI211_X1 g634(.A(G469), .B(new_n303), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n305), .A2(new_n367), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n292), .B2(new_n294), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n720), .A2(new_n672), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n386), .B2(new_n389), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n746), .A2(new_n824), .A3(new_n827), .A4(new_n594), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n818), .B1(new_n828), .B2(new_n787), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n824), .A2(new_n827), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n661), .A3(KEYINPUT42), .A4(new_n814), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT106), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT106), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G131), .ZN(G33));
  NAND3_X1  g651(.A1(new_n830), .A2(new_n661), .A3(new_n733), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G134), .ZN(G36));
  AOI21_X1  g653(.A(new_n672), .B1(new_n386), .B2(new_n389), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n770), .A2(new_n680), .A3(new_n445), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT43), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(KEYINPUT107), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n773), .B1(new_n667), .B2(new_n669), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n848), .B2(KEYINPUT44), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT44), .B2(new_n848), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT45), .B(new_n303), .C1(new_n819), .C2(new_n820), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(G469), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n822), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT46), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n295), .B1(new_n854), .B2(KEYINPUT46), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n308), .B(new_n778), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(G137), .ZN(G39));
  OAI21_X1  g673(.A(new_n308), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  XOR2_X1   g674(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n841), .A2(new_n746), .A3(new_n594), .A4(new_n787), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(G140), .ZN(G42));
  AND2_X1   g680(.A1(new_n846), .A2(new_n472), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n810), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n757), .A2(new_n672), .A3(new_n796), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n305), .B1(new_n292), .B2(KEYINPUT104), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(KEYINPUT104), .B2(new_n292), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n295), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n827), .ZN(new_n878));
  INV_X1    g692(.A(new_n766), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n594), .A3(new_n879), .A4(new_n472), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n470), .A3(new_n680), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n867), .A2(new_n815), .A3(new_n878), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT112), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT112), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT113), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(KEYINPUT113), .ZN(new_n887));
  OAI211_X1 g701(.A(KEYINPUT51), .B(new_n873), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n862), .A2(new_n863), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n877), .A2(new_n720), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n841), .B(new_n868), .C1(new_n891), .C2(KEYINPUT114), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n867), .A2(new_n661), .A3(new_n878), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT48), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n868), .A2(new_n750), .A3(new_n795), .ZN(new_n897));
  OAI211_X1 g711(.A(G952), .B(new_n284), .C1(new_n880), .C2(new_n681), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n885), .A2(new_n873), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n868), .A2(new_n841), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n896), .B(new_n899), .C1(new_n902), .C2(KEYINPUT51), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT115), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n732), .A2(new_n720), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n310), .B1(new_n383), .B2(new_n384), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n387), .B(new_n906), .C1(new_n388), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n696), .A2(new_n706), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n766), .A2(new_n910), .A3(new_n824), .A4(new_n771), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n816), .B(new_n911), .C1(new_n786), .C2(new_n787), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n913), .A2(KEYINPUT52), .A3(new_n754), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT52), .B1(new_n913), .B2(new_n754), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n390), .A2(new_n479), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT110), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n770), .A2(new_n445), .A3(new_n523), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n681), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT110), .B1(new_n470), .B2(new_n680), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n671), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n524), .B(new_n391), .C1(new_n661), .C2(new_n712), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n797), .A2(new_n800), .A3(new_n803), .A4(new_n812), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n830), .A2(new_n814), .A3(new_n815), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n445), .B1(new_n687), .B2(new_n688), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n523), .A3(new_n732), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n752), .A2(new_n746), .A3(new_n840), .A4(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n838), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n834), .A3(new_n835), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n905), .B1(new_n916), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n926), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n911), .A2(KEYINPUT52), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n788), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n754), .A3(new_n816), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n912), .B1(new_n748), .B2(new_n753), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(KEYINPUT52), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n905), .B1(new_n829), .B2(new_n831), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n934), .A2(new_n939), .A3(KEYINPUT111), .A4(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT111), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n913), .A2(new_n754), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT52), .ZN(new_n944));
  INV_X1    g758(.A(new_n816), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n788), .A2(new_n935), .A3(new_n945), .ZN(new_n946));
  AOI22_X1  g760(.A1(new_n943), .A2(new_n944), .B1(new_n946), .B2(new_n754), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n926), .A2(new_n931), .A3(new_n940), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n933), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT54), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n932), .A2(new_n947), .A3(KEYINPUT53), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n916), .A2(new_n932), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(KEYINPUT53), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(KEYINPUT54), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n904), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n894), .A2(new_n903), .A3(KEYINPUT115), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n842), .A2(new_n595), .A3(new_n826), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT109), .Z(new_n960));
  XOR2_X1   g774(.A(new_n876), .B(KEYINPUT49), .Z(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n757), .A3(new_n879), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n348), .A2(new_n365), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n363), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT55), .Z(new_n966));
  XOR2_X1   g780(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n967));
  AND2_X1   g781(.A1(new_n950), .A2(G902), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n966), .B(new_n967), .C1(new_n968), .C2(G210), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n284), .A2(G952), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(G210), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT56), .B1(new_n971), .B2(KEYINPUT116), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(KEYINPUT116), .B2(new_n971), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n969), .B(new_n970), .C1(new_n973), .C2(new_n966), .ZN(G51));
  XNOR2_X1  g788(.A(new_n950), .B(KEYINPUT54), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n822), .B(KEYINPUT57), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n790), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n968), .A2(new_n853), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(G54));
  NAND3_X1  g796(.A1(new_n968), .A2(KEYINPUT58), .A3(G475), .ZN(new_n983));
  INV_X1    g797(.A(new_n465), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT119), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT119), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n970), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(G60));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT59), .Z(new_n991));
  NOR2_X1   g805(.A1(new_n955), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n676), .A2(new_n677), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n991), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n975), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n994), .A2(new_n970), .A3(new_n996), .ZN(G63));
  INV_X1    g811(.A(KEYINPUT122), .ZN(new_n998));
  NAND2_X1  g812(.A1(G217), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT60), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n950), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT120), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n950), .A2(KEYINPUT120), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(KEYINPUT121), .B1(new_n1005), .B2(new_n705), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n950), .A2(KEYINPUT120), .A3(new_n1000), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT120), .B1(new_n950), .B2(new_n1000), .ZN(new_n1008));
  OAI211_X1 g822(.A(KEYINPUT121), .B(new_n705), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n998), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n970), .B1(new_n1012), .B2(new_n590), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT61), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI221_X1 g830(.A(new_n1013), .B1(new_n998), .B2(KEYINPUT61), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G66));
  XNOR2_X1  g832(.A(new_n926), .B(KEYINPUT123), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n352), .A2(new_n284), .ZN(new_n1021));
  AOI22_X1  g835(.A1(new_n1020), .A2(new_n284), .B1(new_n476), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n964), .B1(G898), .B2(new_n284), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(G69));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n284), .A2(G900), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n945), .B(new_n788), .C1(new_n748), .C2(new_n753), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n850), .B2(new_n857), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n857), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1032), .A2(new_n661), .A3(new_n811), .ZN(new_n1033));
  AND4_X1   g847(.A1(new_n836), .A2(new_n865), .A3(new_n838), .A4(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1025), .B(new_n1027), .C1(new_n1035), .C2(G953), .ZN(new_n1036));
  AOI21_X1  g850(.A(G953), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1037));
  OAI21_X1  g851(.A(KEYINPUT126), .B1(new_n1037), .B2(new_n1026), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n626), .B(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1036), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT124), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n784), .A2(new_n1028), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT62), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n780), .A2(new_n662), .A3(new_n841), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1047), .B1(new_n920), .B2(new_n921), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n1046), .A2(new_n858), .A3(new_n865), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n284), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1043), .B1(new_n1050), .B2(new_n1040), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1042), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1052), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1053), .A2(new_n1054), .ZN(G72));
  NAND2_X1  g869(.A1(new_n1035), .A2(new_n1020), .ZN(new_n1056));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT63), .ZN(new_n1058));
  XNOR2_X1  g872(.A(new_n1058), .B(KEYINPUT127), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1060), .A2(new_n644), .A3(new_n742), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1059), .B1(new_n1049), .B2(new_n1019), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(new_n758), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n630), .A2(new_n654), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n1064), .A2(new_n1058), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n970), .B1(new_n954), .B2(new_n1065), .ZN(new_n1066));
  AND3_X1   g880(.A1(new_n1061), .A2(new_n1063), .A3(new_n1066), .ZN(G57));
endmodule


