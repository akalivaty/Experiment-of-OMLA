//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n201), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n211), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n213), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n216), .B(new_n224), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n222), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n204), .A2(new_n211), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n211), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT68), .Z(new_n264));
  NAND3_X1  g0064(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n254), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n267), .B1(new_n202), .B2(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(G223), .B1(new_n280), .B2(G77), .ZN(new_n281));
  INV_X1    g0081(.A(G222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n275), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n272), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n286), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n292), .B(new_n210), .C1(new_n297), .C2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(G226), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n289), .A2(new_n302), .A3(G190), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n269), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n271), .A2(new_n304), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n271), .A4(new_n304), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n303), .A2(G179), .ZN(new_n314));
  AOI21_X1  g0114(.A(G169), .B1(new_n289), .B2(new_n302), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n314), .A2(new_n270), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n277), .A2(G238), .B1(new_n280), .B2(G107), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n238), .B2(new_n284), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n288), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n299), .B1(G244), .B2(new_n301), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n267), .A2(G77), .A3(new_n262), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G77), .B2(new_n265), .ZN(new_n328));
  INV_X1    g0128(.A(new_n258), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n259), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n328), .B1(new_n332), .B2(new_n254), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n324), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n323), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n318), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n275), .A2(new_n211), .A3(new_n276), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT7), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n275), .A2(new_n347), .A3(new_n211), .A4(new_n276), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(G68), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G58), .ZN(new_n350));
  INV_X1    g0150(.A(G68), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n256), .A2(G159), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n353), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n346), .B2(new_n348), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n351), .B1(new_n345), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n359), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n254), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n258), .B1(new_n210), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n267), .B1(new_n266), .B2(new_n258), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n287), .A2(G232), .A3(new_n300), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n287), .A2(new_n300), .A3(KEYINPUT71), .A4(G232), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G87), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n274), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G223), .A2(G1698), .ZN(new_n378));
  INV_X1    g0178(.A(G226), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(G1698), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n283), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n298), .B1(new_n381), .B2(new_n287), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n325), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G223), .B2(G1698), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n280), .B1(new_n274), .B2(new_n376), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n288), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n387), .A2(new_n374), .A3(new_n334), .A4(new_n298), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT72), .B1(new_n369), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n383), .A2(new_n388), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n366), .A3(new_n392), .A4(new_n368), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n344), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n368), .ZN(new_n395));
  INV_X1    g0195(.A(new_n254), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n347), .B1(new_n280), .B2(new_n211), .ZN(new_n397));
  INV_X1    g0197(.A(new_n348), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT70), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n363), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(new_n359), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n395), .B1(new_n401), .B2(new_n358), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n375), .B2(new_n382), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n387), .A2(new_n374), .A3(G179), .A4(new_n298), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT18), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n404), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n369), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT17), .B1(new_n402), .B2(new_n391), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n394), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT67), .B(G41), .ZN(new_n414));
  INV_X1    g0214(.A(G45), .ZN(new_n415));
  AOI21_X1  g0215(.A(G1), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n292), .B1(new_n301), .B2(G238), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n379), .A2(new_n272), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n238), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n278), .C2(new_n279), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n287), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n413), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n287), .A2(G238), .A3(new_n300), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n298), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n426), .A2(KEYINPUT13), .A3(new_n422), .ZN(new_n427));
  OAI21_X1  g0227(.A(G169), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT14), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT13), .B1(new_n426), .B2(new_n422), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT69), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n417), .A2(new_n423), .A3(new_n413), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT69), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(KEYINPUT13), .C1(new_n426), .C2(new_n422), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(G179), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n432), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(G169), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n429), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n351), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n205), .B2(new_n259), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n254), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT11), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n266), .A2(new_n351), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n267), .A2(G68), .A3(new_n262), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n436), .B2(G200), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n431), .A2(G190), .A3(new_n432), .A4(new_n434), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n343), .A2(new_n412), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n210), .B(G45), .C1(new_n458), .C2(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n297), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n288), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(G270), .B1(new_n292), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g0262(.A(G257), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n283), .A2(KEYINPUT75), .A3(G264), .A4(G1698), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT76), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n288), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n469), .ZN(new_n473));
  INV_X1    g0273(.A(new_n465), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n473), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n462), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n477), .B(new_n211), .C1(G33), .C2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  AOI221_X4 g0280(.A(KEYINPUT77), .B1(new_n480), .B2(G20), .C1(new_n253), .C2(new_n222), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT77), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n254), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n479), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT20), .B(new_n479), .C1(new_n481), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n265), .A2(new_n480), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n254), .B(new_n266), .C1(new_n210), .C2(G33), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n480), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n339), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n476), .A2(new_n493), .A3(KEYINPUT21), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n473), .A2(new_n474), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT76), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n470), .A2(new_n471), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n288), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n489), .A2(new_n492), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(G179), .A4(new_n462), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n476), .B2(G200), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n334), .B2(new_n476), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT21), .B1(new_n476), .B2(new_n493), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(KEYINPUT78), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n506), .B(KEYINPUT21), .C1(new_n476), .C2(new_n493), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n501), .B(new_n503), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n211), .B2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n274), .A2(new_n480), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n211), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n211), .A3(G87), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n280), .A2(KEYINPUT22), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n376), .A2(KEYINPUT79), .A3(G20), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n283), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n517), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT24), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n514), .A2(new_n516), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT22), .B1(new_n280), .B2(new_n519), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n283), .A2(new_n521), .A3(new_n522), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT24), .B1(new_n531), .B2(KEYINPUT80), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n524), .A2(new_n525), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n254), .B(new_n527), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT25), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n265), .B2(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n512), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n491), .A2(G107), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n542));
  INV_X1    g0342(.A(G294), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n274), .C2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n461), .A2(G264), .B1(new_n544), .B2(new_n288), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n460), .A2(new_n292), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n339), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n288), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT5), .B1(new_n294), .B2(new_n296), .ZN(new_n549));
  OAI211_X1 g0349(.A(G264), .B(new_n287), .C1(new_n549), .C2(new_n459), .ZN(new_n550));
  AND4_X1   g0350(.A1(G179), .A2(new_n548), .A3(new_n550), .A4(new_n546), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n540), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n550), .A3(new_n546), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G169), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(KEYINPUT81), .C1(new_n337), .C2(new_n553), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n539), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n325), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G190), .B2(new_n553), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n534), .A3(new_n538), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n478), .A2(new_n512), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n207), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n512), .A2(KEYINPUT6), .A3(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n346), .A2(G107), .A3(new_n348), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n254), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n265), .A2(G97), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n491), .B2(G97), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT73), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(new_n287), .C1(new_n549), .C2(new_n459), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n546), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n477), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n288), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n577), .B1(new_n586), .B2(new_n325), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n288), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n546), .A2(new_n578), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(KEYINPUT73), .A3(G200), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(G190), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n576), .A2(new_n587), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n573), .A2(new_n575), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n586), .A2(new_n337), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n339), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n211), .B1(new_n421), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G87), .B2(new_n208), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n259), .B2(new_n478), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n211), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n254), .ZN(new_n605));
  INV_X1    g0405(.A(new_n331), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n267), .B(new_n606), .C1(G1), .C2(new_n274), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n331), .A2(new_n266), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT74), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n604), .A2(new_n254), .B1(new_n266), .B2(new_n331), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT74), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(G250), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n415), .B2(G1), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n210), .A2(new_n290), .A3(G45), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n287), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n277), .A2(G244), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n283), .A2(G238), .A3(new_n272), .ZN(new_n621));
  INV_X1    g0421(.A(new_n515), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n619), .B1(new_n623), .B2(new_n288), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G179), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n339), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n267), .B(G87), .C1(G1), .C2(new_n274), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n605), .A2(new_n608), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n288), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n618), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(G200), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(G190), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n614), .A2(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n598), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n457), .A2(new_n509), .A3(new_n564), .A4(new_n634), .ZN(G372));
  AND3_X1   g0435(.A1(new_n369), .A2(new_n407), .A3(new_n408), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n407), .B1(new_n369), .B2(new_n408), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n392), .B1(new_n402), .B2(new_n391), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n392), .A2(new_n391), .A3(new_n366), .A4(new_n368), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT17), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n411), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n342), .A2(new_n453), .B1(new_n439), .B2(new_n449), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n316), .B1(new_n645), .B2(new_n313), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n609), .A2(new_n610), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT74), .B1(new_n612), .B2(new_n607), .ZN(new_n648));
  AOI211_X1 g0448(.A(new_n337), .B(new_n619), .C1(new_n623), .C2(new_n288), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n339), .B1(new_n629), .B2(new_n618), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n631), .A2(new_n632), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n653), .A2(new_n597), .A3(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT26), .B1(new_n633), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n539), .B1(new_n547), .B2(new_n551), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n501), .B(new_n659), .C1(new_n505), .C2(new_n507), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n593), .A2(new_n633), .A3(new_n559), .A4(new_n597), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n646), .B1(new_n456), .B2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  OAI21_X1  g0467(.A(G213), .B1(new_n667), .B2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT84), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(KEYINPUT84), .A3(KEYINPUT27), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G343), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n539), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n561), .B2(new_n563), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n556), .A2(new_n674), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n665), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n563), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n562), .B1(new_n556), .B2(new_n559), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n679), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(KEYINPUT85), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n675), .A2(new_n499), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n509), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n494), .A2(new_n500), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n476), .A2(new_n493), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n506), .B1(new_n691), .B2(KEYINPUT21), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n504), .A2(KEYINPUT78), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n689), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n694), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n674), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n680), .B2(new_n685), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n659), .A2(new_n675), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n214), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n297), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n220), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT86), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n663), .B2(new_n675), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n661), .B1(new_n694), .B2(new_n659), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT86), .B(new_n674), .C1(new_n715), .C2(new_n658), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT87), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT87), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n713), .A2(new_n719), .A3(new_n714), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n661), .B1(new_n694), .B2(new_n556), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n658), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n723), .A2(new_n714), .A3(new_n675), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT88), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n564), .A2(new_n509), .A3(new_n634), .A4(new_n674), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n586), .A2(new_n649), .A3(new_n545), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  OR3_X1    g0530(.A1(new_n729), .A2(new_n476), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n624), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n476), .A2(new_n553), .A3(new_n590), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n729), .B2(new_n476), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n675), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n727), .B1(new_n728), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n711), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(new_n696), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n211), .A2(G13), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n210), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n706), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G330), .B2(new_n695), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n214), .A2(new_n283), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n214), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n705), .A2(new_n283), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n221), .B2(new_n415), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n248), .A2(new_n415), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n222), .B1(G20), .B2(new_n339), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n748), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n334), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n337), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G97), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G159), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n769), .B1(new_n774), .B2(KEYINPUT32), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT91), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n376), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n775), .B(new_n781), .C1(KEYINPUT32), .C2(new_n774), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n770), .A2(new_n334), .A3(G200), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n211), .A2(new_n337), .A3(KEYINPUT89), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT89), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G20), .B2(G179), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n771), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n283), .B1(new_n512), .B2(new_n783), .C1(new_n789), .C2(new_n205), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n766), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G58), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n782), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n788), .A2(KEYINPUT90), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT90), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n787), .B2(new_n325), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n795), .A2(G190), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n795), .A2(new_n334), .A3(new_n797), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n794), .B1(new_n202), .B2(new_n798), .C1(new_n351), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n798), .B(KEYINPUT92), .ZN(new_n801));
  INV_X1    g0601(.A(G326), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n768), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n543), .B1(new_n783), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n772), .B(KEYINPUT94), .Z(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n791), .ZN(new_n810));
  INV_X1    g0610(.A(new_n789), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n806), .B(new_n810), .C1(G311), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n780), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n283), .B1(new_n813), .B2(G303), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT93), .ZN(new_n815));
  INV_X1    g0615(.A(new_n799), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n814), .A2(KEYINPUT93), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n812), .A2(new_n815), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n800), .B1(new_n803), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n765), .B1(new_n821), .B2(new_n762), .ZN(new_n822));
  INV_X1    g0622(.A(new_n761), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n695), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n750), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  OAI22_X1  g0626(.A1(new_n326), .A2(new_n335), .B1(new_n674), .B2(new_n333), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n341), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n342), .A2(new_n674), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n713), .A2(new_n716), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n341), .A2(new_n675), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n341), .B2(new_n827), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n674), .B(new_n833), .C1(new_n715), .C2(new_n658), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n748), .B1(new_n835), .B2(new_n740), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n831), .A2(new_n739), .A3(new_n834), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n762), .A2(new_n759), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n748), .B1(G77), .B2(new_n840), .C1(new_n833), .C2(new_n760), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n280), .B1(new_n768), .B2(G58), .ZN(new_n842));
  INV_X1    g0642(.A(new_n783), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G68), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n807), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n202), .B2(new_n780), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n798), .B1(new_n799), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT96), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G159), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n853), .B2(new_n791), .C1(new_n854), .C2(new_n789), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n848), .B1(new_n856), .B2(KEYINPUT34), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(KEYINPUT34), .B2(new_n856), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n816), .A2(KEYINPUT95), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n816), .A2(KEYINPUT95), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n805), .ZN(new_n862));
  INV_X1    g0662(.A(G311), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n846), .A2(new_n863), .B1(new_n543), .B2(new_n791), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G116), .B2(new_n811), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n843), .A2(G87), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n769), .A3(new_n280), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n813), .B2(G107), .ZN(new_n868));
  INV_X1    g0668(.A(G303), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n865), .B(new_n868), .C1(new_n869), .C2(new_n798), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n858), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n841), .B1(new_n871), .B2(new_n762), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n838), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n223), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OR3_X1    g0678(.A1(new_n220), .A2(new_n205), .A3(new_n352), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n202), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n210), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n721), .A2(new_n457), .A3(new_n725), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n646), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n673), .A2(G343), .A3(new_n449), .ZN(new_n885));
  AOI221_X4 g0685(.A(new_n885), .B1(new_n451), .B2(new_n452), .C1(new_n439), .C2(new_n449), .ZN(new_n886));
  INV_X1    g0686(.A(new_n885), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n450), .B2(new_n453), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n660), .A2(new_n662), .ZN(new_n891));
  INV_X1    g0691(.A(new_n651), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n654), .B1(new_n653), .B2(new_n597), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n633), .A2(new_n656), .A3(KEYINPUT26), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n675), .B(new_n830), .C1(new_n891), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n829), .B(KEYINPUT97), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n890), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n639), .A2(new_n640), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n400), .B2(new_n355), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n365), .A2(new_n254), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n368), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT98), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT98), .B(new_n368), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n408), .C2(new_n673), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n390), .A2(new_n393), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n369), .A2(new_n408), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n369), .A2(new_n673), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n909), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n641), .A2(new_n638), .A3(new_n642), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n905), .A2(new_n673), .A3(new_n906), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n916), .A2(KEYINPUT99), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT99), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  OAI211_X1 g0720(.A(KEYINPUT38), .B(new_n915), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n899), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n638), .A2(new_n673), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT100), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n921), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n916), .A2(new_n369), .A3(new_n673), .ZN(new_n929));
  INV_X1    g0729(.A(new_n914), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT101), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n900), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT101), .B1(new_n910), .B2(new_n914), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n911), .B(new_n912), .C1(new_n369), .C2(new_n389), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT37), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n923), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n921), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n450), .A2(new_n675), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n928), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n889), .B1(new_n834), .B2(new_n897), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT99), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n412), .B2(new_n917), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n916), .A2(KEYINPUT99), .A3(new_n918), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n948), .B2(new_n915), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n908), .A2(KEYINPUT37), .B1(new_n900), .B2(new_n930), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n923), .B(new_n950), .C1(new_n946), .C2(new_n947), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n944), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT100), .ZN(new_n953));
  INV_X1    g0753(.A(new_n926), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n927), .A2(new_n943), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n884), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n833), .B1(new_n886), .B2(new_n888), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n728), .B2(new_n738), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n949), .B2(new_n951), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n929), .B2(new_n936), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n950), .B1(new_n946), .B2(new_n947), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(KEYINPUT38), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(KEYINPUT40), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n728), .A2(new_n738), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n457), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(G330), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n957), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n210), .B2(new_n745), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n957), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n882), .B1(new_n974), .B2(new_n975), .ZN(G367));
  OAI21_X1  g0776(.A(new_n598), .B1(new_n576), .B2(new_n674), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n656), .A2(new_n675), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n701), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT42), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n597), .B1(new_n977), .B2(new_n556), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT102), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n674), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n980), .B2(KEYINPUT42), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n675), .A2(new_n628), .ZN(new_n987));
  MUX2_X1   g0787(.A(new_n892), .B(new_n633), .S(new_n987), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n981), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n697), .A2(new_n979), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n989), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n993), .B1(new_n991), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n706), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(new_n979), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n701), .B2(new_n702), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n700), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n686), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n702), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n1005), .A3(new_n979), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT103), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT103), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n703), .A2(new_n1008), .A3(new_n979), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1009), .A3(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT45), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n697), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1012), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1014), .A2(new_n698), .A3(new_n1002), .A4(new_n1010), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n687), .A2(new_n700), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n744), .A3(new_n1004), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n686), .A2(new_n1003), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n696), .B1(new_n1018), .B2(new_n701), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n741), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1013), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n998), .B1(new_n1022), .B2(new_n742), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n997), .B1(new_n1023), .B2(new_n747), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n813), .A2(G116), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT46), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT104), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G283), .A2(new_n811), .B1(new_n792), .B2(G303), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n280), .B1(new_n772), .B2(new_n1030), .C1(new_n478), .C2(new_n783), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G107), .B2(new_n768), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(new_n1026), .C2(new_n1025), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n863), .B2(new_n801), .C1(new_n861), .C2(new_n543), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n280), .B1(new_n773), .B2(G137), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n205), .B2(new_n783), .C1(new_n351), .C2(new_n804), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n202), .A2(new_n789), .B1(new_n791), .B2(new_n850), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G58), .C2(new_n813), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n853), .B2(new_n801), .C1(new_n861), .C2(new_n854), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT47), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT47), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n762), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n748), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n754), .A2(new_n244), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n764), .B1(new_n705), .B2(new_n606), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1044), .B(new_n1048), .C1(new_n823), .C2(new_n988), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1024), .A2(new_n1049), .ZN(G387));
  NOR2_X1   g0850(.A1(new_n1020), .A2(new_n746), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT105), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n687), .A2(new_n761), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n751), .A2(new_n708), .B1(G107), .B2(new_n214), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n241), .A2(new_n415), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n708), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n1056), .C1(G68), .C2(G77), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n258), .A2(G50), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n755), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1054), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n748), .B1(new_n1061), .B2(new_n764), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n799), .A2(new_n258), .B1(new_n351), .B2(new_n789), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT107), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n768), .A2(new_n606), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n791), .B2(new_n202), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT106), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n813), .A2(G77), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n280), .B1(new_n773), .B2(G150), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n478), .C2(new_n783), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n798), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(G159), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1064), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n283), .B1(new_n773), .B2(G326), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n780), .A2(new_n543), .B1(new_n805), .B2(new_n804), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT108), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n869), .A2(new_n789), .B1(new_n791), .B2(new_n1030), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT109), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n809), .B2(new_n801), .C1(new_n861), .C2(new_n863), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT48), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT49), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1074), .B1(new_n480), .B2(new_n783), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1073), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1062), .B1(new_n1086), .B2(new_n762), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1052), .B1(new_n1053), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1021), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n741), .A2(new_n1020), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n706), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(G393));
  NAND3_X1  g0892(.A1(new_n1013), .A2(new_n1015), .A3(new_n747), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n789), .A2(new_n543), .B1(new_n480), .B2(new_n804), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n283), .B1(new_n773), .B2(G322), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n512), .B2(new_n783), .C1(new_n780), .C2(new_n805), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT112), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n798), .A2(new_n1030), .B1(new_n863), .B2(new_n791), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1099));
  AOI211_X1 g0899(.A(new_n1094), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n869), .B2(new_n861), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT113), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n798), .A2(new_n850), .B1(new_n854), .B2(new_n791), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT51), .Z(new_n1104));
  AOI21_X1  g0904(.A(new_n280), .B1(new_n773), .B2(G143), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n768), .A2(G77), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n866), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n789), .A2(new_n258), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G68), .C2(new_n813), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n861), .B2(new_n202), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1102), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1101), .A2(KEYINPUT113), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n762), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n754), .A2(new_n251), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1114), .B(new_n763), .C1(new_n478), .C2(new_n214), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT110), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1117), .A2(new_n1118), .A3(new_n1045), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1113), .B(new_n1119), .C1(new_n823), .C2(new_n979), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1022), .A2(new_n706), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1021), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1093), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(G390));
  NAND3_X1  g0923(.A1(new_n739), .A2(new_n833), .A3(new_n890), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n674), .B(new_n828), .C1(new_n722), .C2(new_n658), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n889), .B1(new_n1125), .B2(new_n829), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n965), .A2(new_n1126), .A3(new_n942), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n928), .A2(new_n941), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n834), .A2(new_n897), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n942), .B1(new_n1130), .B2(new_n890), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1124), .B(new_n1128), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1124), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n928), .B2(new_n941), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n747), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1045), .B1(new_n258), .B2(new_n839), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n861), .A2(new_n849), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n780), .A2(new_n850), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1071), .A2(G128), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n847), .A2(new_n791), .B1(new_n789), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G125), .B2(new_n807), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n283), .B1(new_n804), .B2(new_n854), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G50), .B2(new_n843), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n861), .A2(new_n512), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n478), .A2(new_n789), .B1(new_n791), .B2(new_n480), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G294), .B2(new_n807), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n844), .A2(new_n1106), .A3(new_n280), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n781), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n805), .C2(new_n798), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1138), .A2(new_n1147), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n762), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1137), .B1(new_n1155), .B2(new_n1157), .C1(new_n1129), .C2(new_n760), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1136), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT116), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1136), .A2(KEYINPUT116), .A3(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n890), .B1(new_n739), .B2(new_n833), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1130), .B1(new_n1133), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1125), .A2(new_n829), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1124), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n457), .A2(new_n739), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1169), .A2(new_n883), .A3(new_n646), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n706), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT114), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT114), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n706), .C1(new_n1163), .C2(new_n1171), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1163), .A2(new_n1171), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1161), .B(new_n1162), .C1(new_n1174), .C2(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(new_n673), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n270), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n318), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT119), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1181), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n313), .A2(new_n317), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n313), .B2(new_n317), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1181), .B(new_n316), .C1(new_n309), .C2(new_n312), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT119), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1190));
  AND3_X1   g0990(.A1(new_n1186), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n924), .A2(new_n921), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT40), .B1(new_n1195), .B2(new_n959), .ZN(new_n1196));
  OAI21_X1  g0996(.A(G330), .B1(new_n965), .B2(new_n966), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n961), .B(new_n958), .C1(new_n728), .C2(new_n738), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n727), .B1(new_n939), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n958), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n968), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n924), .B2(new_n921), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n1193), .C1(new_n1203), .C2(KEYINPUT40), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(new_n956), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n955), .A2(new_n943), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(new_n927), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n883), .A2(new_n646), .A3(new_n1170), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1169), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n706), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1205), .A2(new_n956), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT120), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT121), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1204), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1193), .B1(new_n962), .B2(new_n1200), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1207), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1218), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1205), .A2(new_n956), .A3(KEYINPUT121), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1217), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1211), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1169), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1163), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT121), .B1(new_n1205), .B2(new_n956), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1223), .A2(new_n1218), .A3(new_n1204), .A4(new_n1198), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT120), .B1(new_n1205), .B2(new_n956), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1226), .A2(new_n1229), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1214), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1226), .A2(new_n747), .A3(new_n1233), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1194), .A2(new_n759), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n283), .A2(new_n297), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1068), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT118), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1240), .A2(new_n1241), .B1(G97), .B2(new_n816), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n480), .B2(new_n798), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G107), .A2(new_n792), .B1(new_n811), .B2(new_n606), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G58), .A2(new_n843), .B1(new_n768), .B2(G68), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n805), .C2(new_n846), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1243), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT58), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G50), .B(new_n1239), .C1(new_n274), .C2(new_n293), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT117), .Z(new_n1251));
  AND2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n780), .A2(new_n1142), .ZN(new_n1253));
  INV_X1    g1053(.A(G128), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n791), .A2(new_n1254), .B1(new_n850), .B2(new_n804), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1253), .B(new_n1255), .C1(G137), .C2(new_n811), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1071), .A2(G125), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n847), .C2(new_n799), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n843), .A2(G159), .ZN(new_n1261));
  AOI211_X1 g1061(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1252), .B1(KEYINPUT58), .B2(new_n1248), .C1(new_n1259), .C2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n762), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n839), .A2(new_n202), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1238), .A2(new_n748), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1237), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1236), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(G375));
  NAND2_X1  g1070(.A1(new_n1211), .A2(new_n1228), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT122), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n998), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT122), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1211), .A2(new_n1274), .A3(new_n1228), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1171), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1169), .A2(new_n747), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n748), .B1(G68), .B2(new_n840), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT123), .Z(new_n1279));
  AOI22_X1  g1079(.A1(new_n1071), .A2(G294), .B1(G107), .B2(new_n811), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n861), .B2(new_n480), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT124), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1065), .B(new_n280), .C1(new_n205), .C2(new_n783), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n846), .A2(new_n869), .B1(new_n805), .B2(new_n791), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(G97), .C2(new_n813), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n846), .A2(new_n1254), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n849), .A2(new_n791), .B1(new_n789), .B2(new_n850), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n780), .A2(new_n854), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n283), .B1(new_n783), .B2(new_n350), .C1(new_n804), .C2(new_n202), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n847), .B2(new_n798), .C1(new_n861), .C2(new_n1142), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n762), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1279), .B1(new_n760), .B2(new_n890), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1276), .A2(new_n1297), .ZN(G381));
  NAND3_X1  g1098(.A1(new_n1088), .A2(new_n825), .A3(new_n1091), .ZN(new_n1299));
  OR4_X1    g1099(.A1(G384), .A2(G390), .A3(new_n1299), .A4(G381), .ZN(new_n1300));
  OR3_X1    g1100(.A1(new_n1300), .A2(KEYINPUT125), .A3(G387), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT125), .B1(new_n1300), .B2(G387), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1136), .B(new_n1158), .C1(new_n1174), .C2(new_n1178), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1301), .A2(new_n1269), .A3(new_n1302), .A4(new_n1304), .ZN(G407));
  NAND2_X1  g1105(.A1(new_n1269), .A2(new_n1304), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G343), .C2(new_n1306), .ZN(G409));
  INV_X1    g1107(.A(G343), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(G213), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1272), .A2(new_n1275), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1271), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n707), .B1(new_n1312), .B2(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1314), .B2(new_n1297), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n873), .B(new_n1296), .C1(new_n1311), .C2(new_n1313), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1173), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1236), .A2(new_n1268), .A3(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1267), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1323), .B2(new_n1215), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(new_n746), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(KEYINPUT126), .A3(new_n1215), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1322), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1226), .A2(new_n1229), .A3(new_n1233), .A4(new_n1273), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1303), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1309), .B(new_n1317), .C1(new_n1321), .C2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1309), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1314), .A2(new_n1297), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n873), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1314), .A2(G384), .A3(new_n1297), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1308), .A2(G213), .A3(G2897), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1336), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1332), .A2(new_n1340), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1232), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1322), .B1(new_n1344), .B2(new_n747), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT57), .B1(new_n1344), .B2(new_n1229), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G378), .B(new_n1345), .C1(new_n1346), .C2(new_n1214), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1304), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1350), .A2(new_n1351), .A3(new_n1309), .A4(new_n1317), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT61), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1331), .A2(new_n1341), .A3(new_n1352), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G393), .A2(G396), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1299), .ZN(new_n1356));
  AND3_X1   g1156(.A1(new_n1024), .A2(new_n1049), .A3(G390), .ZN(new_n1357));
  AOI21_X1  g1157(.A(G390), .B1(new_n1024), .B2(new_n1049), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1356), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(G390), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G387), .A2(new_n1360), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1355), .A2(new_n1299), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1024), .A2(new_n1049), .A3(G390), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1359), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1354), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT63), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1365), .B1(new_n1367), .B2(new_n1330), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1330), .A2(new_n1367), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT61), .B1(new_n1332), .B2(new_n1340), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1368), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1366), .A2(new_n1371), .ZN(G405));
  INV_X1    g1172(.A(new_n1317), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1365), .A2(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1359), .A2(new_n1364), .A3(new_n1317), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1304), .B1(new_n1236), .B2(new_n1268), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1347), .A2(new_n1376), .A3(KEYINPUT127), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1377), .B1(KEYINPUT127), .B2(new_n1376), .ZN(new_n1378));
  AND3_X1   g1178(.A1(new_n1374), .A2(new_n1375), .A3(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1378), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1380));
  NOR2_X1   g1180(.A1(new_n1379), .A2(new_n1380), .ZN(G402));
endmodule


