//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(KEYINPUT68), .A3(G101), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n469), .A2(G137), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(G160));
  NAND2_X1  g053(.A1(new_n469), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT70), .B1(new_n468), .B2(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n462), .A2(new_n484), .A3(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(G124), .B2(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT71), .B1(new_n462), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(KEYINPUT71), .B(new_n492), .C1(new_n466), .C2(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n462), .A2(G138), .A3(new_n464), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n462), .A2(new_n501), .A3(G138), .A4(new_n464), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(KEYINPUT72), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n508), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n515), .A2(G88), .B1(G50), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(new_n523), .A3(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  OAI211_X1 g100(.A(G50), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n519), .B1(new_n513), .B2(new_n512), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n529), .B2(new_n522), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(new_n514), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n511), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n537), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  OAI211_X1 g118(.A(G52), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n509), .B2(new_n510), .ZN(new_n548));
  AND2_X1   g123(.A1(G77), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n543), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n515), .A2(G90), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n553), .A2(KEYINPUT74), .A3(new_n550), .A4(new_n544), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(G171));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G43), .Z(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n535), .A2(new_n556), .B1(new_n527), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n518), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  AOI22_X1  g141(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n518), .ZN(new_n568));
  OAI211_X1 g143(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n515), .A2(G91), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT76), .A4(new_n571), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  NAND3_X1  g154(.A1(new_n524), .A2(new_n530), .A3(KEYINPUT77), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT77), .B1(new_n524), .B2(new_n530), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n515), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n516), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n519), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(G73), .A3(G543), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n518), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n509), .B2(new_n510), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n592), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n595), .B(G651), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n534), .A2(G86), .A3(new_n519), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n534), .A2(G48), .A3(G543), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n596), .A2(new_n603), .ZN(G305));
  XNOR2_X1  g179(.A(KEYINPUT80), .B(G47), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n535), .A2(new_n605), .B1(new_n527), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n518), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(new_n516), .A2(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n518), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n527), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n620), .B(G301), .S(G868), .Z(G284));
  XOR2_X1   g196(.A(G284), .B(KEYINPUT81), .Z(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n619), .A2(new_n627), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT82), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(KEYINPUT83), .C1(G868), .C2(new_n561), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(KEYINPUT83), .B2(new_n631), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n462), .A2(new_n471), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n469), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n464), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G123), .B2(new_n486), .ZN(new_n645));
  AOI22_X1  g220(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n640), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n647), .C1(new_n639), .C2(new_n638), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n661), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n639), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n640), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT86), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G5), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G171), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1961), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  INV_X1    g276(.A(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n702), .B2(KEYINPUT24), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(KEYINPUT24), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G160), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n699), .B2(G1961), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT25), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n469), .A2(G139), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n464), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n706), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n706), .B2(G33), .ZN(new_n719));
  INV_X1    g294(.A(G2072), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n697), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n697), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G1966), .ZN(new_n724));
  INV_X1    g299(.A(G11), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT31), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G28), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n706), .B1(new_n728), .B2(G28), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n727), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n645), .B2(G29), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n721), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n707), .A2(new_n708), .ZN(new_n734));
  OR4_X1    g309(.A1(new_n701), .A2(new_n710), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n719), .A2(new_n720), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n706), .A2(G32), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n486), .A2(G129), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n469), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n471), .A2(G105), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(new_n706), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n723), .A2(G1966), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT92), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n706), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n706), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n737), .A2(new_n748), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n735), .A2(new_n755), .A3(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n697), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n624), .B2(new_n697), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1956), .Z(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G162), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n619), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G4), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n706), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n486), .A2(G128), .ZN(new_n772));
  NOR2_X1   g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT89), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n470), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G140), .ZN(new_n778));
  INV_X1    g353(.A(new_n469), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n772), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n771), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n767), .A2(new_n768), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n697), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n561), .B2(new_n697), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n769), .A2(new_n783), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n760), .A2(new_n765), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n756), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G22), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G166), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(G6), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G305), .B2(new_n697), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n697), .A2(G23), .ZN(new_n801));
  INV_X1    g376(.A(G288), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n697), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT88), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n794), .A2(new_n799), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n809));
  NOR2_X1   g384(.A1(G25), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n486), .A2(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT87), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n470), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI22_X1  g390(.A1(G131), .A2(new_n469), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(G29), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n697), .A2(G24), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n610), .B2(new_n697), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n809), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT94), .B1(new_n735), .B2(new_n755), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n790), .A2(new_n829), .A3(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  AOI22_X1  g407(.A1(new_n515), .A2(G93), .B1(G55), .B2(new_n516), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT95), .B1(new_n834), .B2(new_n518), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n834), .A2(KEYINPUT95), .A3(new_n518), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n561), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n558), .B2(new_n560), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n836), .A2(new_n839), .A3(new_n561), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT38), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n627), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n838), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n645), .B(KEYINPUT97), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n705), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n469), .A2(G142), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n486), .A2(G130), .ZN(new_n860));
  OR2_X1    g435(.A1(G106), .A2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(new_n637), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n859), .A2(new_n866), .A3(new_n860), .A4(new_n862), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n865), .B1(new_n864), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n817), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n818), .A3(new_n868), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n745), .B(new_n780), .ZN(new_n874));
  INV_X1    g449(.A(new_n717), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n492), .B1(new_n466), .B2(new_n467), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT71), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n490), .B1(new_n879), .B2(new_n494), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n880), .A2(new_n881), .B1(new_n500), .B2(new_n502), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n496), .A2(KEYINPUT98), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI22_X1  g460(.A1(G140), .A2(new_n469), .B1(new_n774), .B2(new_n776), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n745), .A2(new_n772), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n780), .B1(new_n739), .B2(new_n744), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n717), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n876), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n885), .B1(new_n876), .B2(new_n890), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n871), .B(new_n873), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n876), .A2(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n884), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n891), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(KEYINPUT101), .A3(new_n873), .A4(new_n871), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n871), .A2(new_n873), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n891), .A3(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n896), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n856), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n899), .A2(KEYINPUT103), .B1(new_n873), .B2(new_n871), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n856), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n896), .A2(new_n900), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT40), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G395));
  NOR2_X1   g490(.A1(G166), .A2(new_n802), .ZN(new_n916));
  AOI21_X1  g491(.A(G288), .B1(new_n524), .B2(new_n530), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G305), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n922), .A2(KEYINPUT107), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(KEYINPUT42), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT107), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n844), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n630), .B(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n574), .A2(new_n576), .A3(new_n619), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n619), .B1(new_n574), .B2(new_n576), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  INV_X1    g512(.A(new_n932), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n930), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(new_n933), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n929), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n927), .B(new_n945), .ZN(new_n946));
  MUX2_X1   g521(.A(new_n838), .B(new_n946), .S(G868), .Z(G295));
  MUX2_X1   g522(.A(new_n838), .B(new_n946), .S(G868), .Z(G331));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n552), .A2(new_n554), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G286), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n953), .A3(G286), .ZN(new_n954));
  NAND2_X1  g529(.A1(G171), .A2(KEYINPUT108), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n844), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n950), .A2(new_n953), .A3(G286), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n953), .B1(new_n950), .B2(G286), .ZN(new_n960));
  OAI211_X1 g535(.A(G171), .B(KEYINPUT108), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n928), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n933), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n939), .B1(new_n938), .B2(new_n930), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n936), .B2(new_n933), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n958), .A3(new_n963), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n967), .A2(new_n958), .A3(KEYINPUT110), .A4(new_n963), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n922), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n958), .B(new_n963), .C1(new_n942), .C2(new_n943), .ZN(new_n972));
  INV_X1    g547(.A(new_n933), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n961), .A2(new_n928), .A3(new_n962), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n928), .B1(new_n961), .B2(new_n962), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n976), .A3(new_n922), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT111), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n968), .A2(new_n965), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n976), .A3(new_n970), .ZN(new_n982));
  INV_X1    g557(.A(new_n922), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n977), .A2(new_n978), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n987), .A3(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n922), .B1(new_n972), .B2(new_n976), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n979), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n984), .A2(new_n985), .A3(new_n992), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n992), .B2(new_n991), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n989), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(G397));
  XOR2_X1   g573(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n881), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n503), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n880), .A2(new_n881), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n465), .A2(new_n476), .A3(G40), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n745), .B(G1996), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n780), .B(new_n782), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n818), .A2(new_n821), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n818), .A2(new_n821), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1986), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n610), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n882), .B2(new_n883), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1009), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT115), .B(G8), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n802), .A2(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n596), .A2(new_n603), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n594), .A2(new_n595), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n1030));
  OAI21_X1  g605(.A(G1981), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(new_n1031), .A3(KEYINPUT49), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(new_n1023), .A3(new_n1021), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1026), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1026), .A2(new_n1036), .A3(KEYINPUT118), .A4(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT45), .B(new_n1001), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n880), .A2(KEYINPUT72), .B1(new_n500), .B2(new_n502), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n1046), .B2(new_n498), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n1020), .C1(new_n1047), .C2(new_n1000), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n793), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1009), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n504), .A2(new_n503), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n880), .A2(KEYINPUT72), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1052), .B(new_n1001), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1053), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1049), .B1(new_n1058), .B2(G2090), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1023), .ZN(new_n1060));
  NAND4_X1  g635(.A1(G303), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT77), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G166), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(G8), .A3(new_n580), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1060), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1020), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n764), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1075), .B2(new_n1049), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1069), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT45), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1005), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n505), .A2(new_n1001), .A3(new_n1000), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1020), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1966), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1009), .B1(new_n1019), .B2(new_n1052), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n505), .A2(new_n1001), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT50), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1087), .A3(new_n708), .ZN(new_n1088));
  AOI211_X1 g663(.A(G286), .B(new_n1022), .C1(new_n1084), .C2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1044), .A2(new_n1070), .A3(new_n1078), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1040), .A2(new_n1091), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n1078), .A3(new_n1089), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1021), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(new_n1022), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1036), .A2(new_n1037), .A3(new_n802), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1028), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1078), .B2(new_n1040), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1100), .B(new_n1103), .C1(new_n1078), .C2(new_n1040), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1092), .A2(new_n1095), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT119), .B(G1956), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1058), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1009), .B1(new_n1019), .B2(KEYINPUT45), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1108), .B(new_n1109), .C1(new_n1047), .C2(new_n1000), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n572), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT57), .A4(new_n571), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n572), .A2(KEYINPUT121), .A3(new_n1111), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1107), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1048), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1058), .A2(new_n1106), .B1(new_n1119), .B2(new_n1109), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1114), .A2(new_n1115), .A3(KEYINPUT123), .A4(new_n1116), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n1131));
  AOI21_X1  g706(.A(G1348), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1021), .A2(G2067), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1096), .A2(new_n782), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(KEYINPUT122), .C1(new_n1074), .C2(G1348), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1136), .A3(new_n619), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1118), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1117), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1118), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT58), .B(G1341), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1048), .A2(G1996), .B1(new_n1096), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n561), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1146), .A3(new_n561), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1107), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT61), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n620), .B1(new_n1154), .B2(KEYINPUT60), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1156), .B(new_n619), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1155), .A2(new_n1157), .B1(KEYINPUT60), .B2(new_n1154), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1138), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT125), .B(KEYINPUT51), .Z(new_n1160));
  AOI21_X1  g735(.A(new_n1071), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G286), .A2(new_n1023), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1160), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT126), .B(new_n1160), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n1023), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1166), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1170), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1162), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1042), .A2(new_n1043), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT53), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1048), .B2(G2078), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1074), .A2(G1961), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g758(.A(G171), .B(KEYINPUT54), .Z(new_n1184));
  NOR2_X1   g759(.A1(new_n1179), .A2(G2078), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1108), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1186), .B2(new_n1008), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1080), .A2(new_n1081), .A3(new_n1020), .A4(new_n1185), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1180), .B(new_n1188), .C1(new_n1074), .C2(G1961), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1183), .A2(new_n1187), .B1(new_n1189), .B2(new_n1184), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1178), .A2(new_n1190), .A3(new_n1070), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1105), .B1(new_n1159), .B2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1189), .A2(G171), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1178), .A2(new_n1070), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1171), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1175), .B1(new_n1196), .B2(new_n1167), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g774(.A(KEYINPUT62), .B(new_n1175), .C1(new_n1196), .C2(new_n1167), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1018), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1012), .A2(new_n745), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1010), .A2(new_n1203), .ZN(new_n1204));
  OR3_X1    g779(.A1(new_n1008), .A2(G1996), .A3(new_n1009), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1205), .A2(KEYINPUT46), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(KEYINPUT46), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT47), .Z(new_n1209));
  XOR2_X1   g784(.A(new_n1013), .B(KEYINPUT127), .Z(new_n1210));
  NAND2_X1  g785(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1211));
  OAI22_X1  g786(.A1(new_n1210), .A2(new_n1211), .B1(G2067), .B2(new_n780), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1212), .A2(new_n1010), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1010), .A2(new_n1016), .A3(new_n610), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT48), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1217), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1213), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1209), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1202), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g796(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n695), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n907), .B2(new_n912), .ZN(new_n1225));
  AND2_X1   g799(.A1(new_n1225), .A2(new_n996), .ZN(G308));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n996), .ZN(G225));
endmodule


