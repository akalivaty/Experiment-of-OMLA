//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT70), .Z(G217));
  OR4_X1    g029(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT71), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  NAND2_X1  g036(.A1(new_n456), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT72), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n470), .B1(new_n473), .B2(KEYINPUT73), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G125), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g052(.A(G137), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n482), .ZN(G160));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n479), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n468), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n471), .A2(new_n472), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(G136), .B2(new_n493), .ZN(G162));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT74), .A2(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n468), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT3), .B(G2104), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G138), .A4(new_n468), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n504), .B2(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  AND3_X1   g094(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n518), .A2(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n516), .A2(new_n526), .ZN(G166));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n510), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n511), .A2(new_n512), .B1(new_n528), .B2(new_n529), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n515), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(G90), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n518), .A2(new_n541), .B1(new_n524), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n515), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT77), .B(G43), .Z(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n518), .A2(new_n547), .B1(new_n524), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n520), .A2(new_n521), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n513), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n518), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n530), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n567), .B1(G91), .B2(new_n536), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT79), .Z(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n511), .A2(new_n574), .A3(new_n512), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n536), .A2(G87), .B1(new_n575), .B2(G651), .ZN(new_n576));
  OAI211_X1 g151(.A(G49), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n517), .A2(KEYINPUT80), .A3(G49), .A4(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G288));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n557), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n513), .A2(KEYINPUT81), .A3(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n518), .A2(new_n590), .B1(new_n524), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n515), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n518), .A2(new_n597), .B1(new_n524), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n530), .A2(G54), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n536), .B2(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n558), .A2(new_n560), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT82), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n515), .B1(new_n608), .B2(KEYINPUT82), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n569), .B(KEYINPUT79), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n487), .A2(G123), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT83), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n493), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n468), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT84), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n505), .A2(new_n480), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n643));
  OAI22_X1  g218(.A1(new_n642), .A2(new_n643), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n650), .A2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT89), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n675), .A2(new_n680), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n690), .B2(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(G127), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n492), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g273(.A1(G115), .A2(G2104), .ZN(new_n699));
  OAI21_X1  g274(.A(G2105), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT94), .B(KEYINPUT25), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n493), .A2(G139), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G33), .ZN(new_n710));
  INV_X1    g285(.A(G2072), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(G32), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G129), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n480), .A2(G105), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n505), .A2(new_n468), .ZN(new_n719));
  INV_X1    g294(.A(G141), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n713), .B1(new_n722), .B2(new_n709), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n629), .A2(new_n709), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n709), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n712), .A2(new_n725), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT98), .B(G1966), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n709), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G160), .B2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT97), .B(G2084), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n736), .B(new_n743), .C1(new_n710), .C2(new_n711), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n732), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n732), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G1961), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT99), .Z(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G35), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G162), .B2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT29), .B(G2090), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G27), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n756), .C1(G1961), .C2(new_n746), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n731), .A2(new_n744), .A3(new_n748), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n732), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT23), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1956), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n611), .A2(G16), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G4), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1348), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n732), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n550), .B2(new_n732), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1341), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n709), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n493), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n487), .A2(G128), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n772), .B1(new_n778), .B2(new_n709), .ZN(new_n779));
  INV_X1    g354(.A(G2067), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n766), .A2(new_n767), .A3(new_n770), .A4(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n758), .B(new_n762), .C1(new_n782), .C2(KEYINPUT93), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(KEYINPUT93), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n732), .A2(G24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n600), .B2(new_n732), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1986), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n487), .A2(G119), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n468), .A2(G107), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n790));
  INV_X1    g365(.A(G131), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n788), .B1(new_n789), .B2(new_n790), .C1(new_n791), .C2(new_n719), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n787), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n732), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n732), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n732), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n732), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(new_n801), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n797), .B1(new_n796), .B2(new_n794), .C1(new_n811), .C2(KEYINPUT34), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(KEYINPUT34), .B2(new_n811), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT36), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n784), .A2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  XNOR2_X1  g391(.A(KEYINPUT101), .B(G860), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n611), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(G80), .A2(G543), .ZN(new_n821));
  INV_X1    g396(.A(G67), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n557), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(new_n821), .C1(new_n557), .C2(new_n822), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n826), .A3(G651), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n536), .A2(G93), .B1(new_n530), .B2(G55), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n550), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n820), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n818), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(new_n818), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n792), .B(new_n633), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n487), .A2(G130), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT102), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G118), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n493), .B2(G142), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n839), .A2(new_n841), .A3(new_n845), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(KEYINPUT103), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT103), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n504), .A2(new_n507), .ZN(new_n852));
  AND2_X1   g427(.A1(KEYINPUT74), .A2(G114), .ZN(new_n853));
  NOR2_X1   g428(.A1(KEYINPUT74), .A2(G114), .ZN(new_n854));
  OAI21_X1  g429(.A(G2105), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n501), .ZN(new_n856));
  AOI22_X1  g431(.A1(G126), .A2(new_n487), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n777), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n707), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n722), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n722), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n851), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n860), .A2(new_n722), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n865), .A2(new_n861), .A3(new_n848), .A4(new_n847), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n629), .B(G160), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(G162), .Z(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT104), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n865), .B(new_n861), .C1(new_n849), .C2(new_n850), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n868), .B1(new_n874), .B2(new_n864), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(G37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT40), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(G166), .B(KEYINPUT107), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(new_n807), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n807), .ZN(new_n886));
  XNOR2_X1  g461(.A(G305), .B(new_n600), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(KEYINPUT108), .A3(new_n889), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT108), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(KEYINPUT42), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n620), .B(new_n831), .ZN(new_n897));
  INV_X1    g472(.A(new_n611), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n615), .ZN(new_n900));
  NAND2_X1  g475(.A1(G299), .A2(KEYINPUT106), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(G299), .A2(KEYINPUT106), .A3(new_n898), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n897), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n896), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n896), .B1(new_n904), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n829), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(G868), .B2(new_n914), .ZN(G295));
  OAI21_X1  g490(.A(new_n913), .B1(G868), .B2(new_n914), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NOR2_X1   g492(.A1(G168), .A2(KEYINPUT109), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n831), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n831), .A2(new_n918), .ZN(new_n920));
  AOI21_X1  g495(.A(G301), .B1(KEYINPUT109), .B2(G168), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n907), .A2(new_n925), .A3(new_n909), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n903), .A4(new_n902), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n928), .B2(new_n895), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n894), .A3(new_n927), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n917), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT54), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT110), .B(G40), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n478), .A2(new_n481), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n477), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G125), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n485), .B2(new_n486), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n469), .B1(new_n946), .B2(new_n475), .ZN(new_n947));
  INV_X1    g522(.A(new_n476), .ZN(new_n948));
  OAI21_X1  g523(.A(G2105), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n943), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT111), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n852), .B2(new_n857), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n944), .A2(new_n951), .B1(KEYINPUT45), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT113), .B(new_n954), .C1(G164), .C2(G1384), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n952), .B2(KEYINPUT45), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n953), .A2(new_n755), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n960));
  AOI211_X1 g535(.A(G1384), .B(new_n960), .C1(new_n852), .C2(new_n857), .ZN(new_n961));
  INV_X1    g536(.A(new_n952), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(KEYINPUT50), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n944), .A2(new_n951), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1961), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n958), .A2(new_n959), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT124), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT111), .B1(new_n949), .B2(new_n950), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n476), .A3(new_n469), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n941), .B(new_n943), .C1(new_n973), .C2(G2105), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n975), .B2(G2078), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n858), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n954), .B(G1384), .C1(new_n852), .C2(new_n857), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(KEYINPUT124), .A3(new_n755), .A4(new_n964), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(KEYINPUT53), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G301), .B1(new_n967), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n958), .A2(new_n959), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n755), .A2(KEYINPUT53), .A3(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n477), .A2(new_n482), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n980), .A2(KEYINPUT125), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n969), .A2(new_n970), .A3(new_n986), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n965), .A2(new_n966), .ZN(new_n992));
  AND4_X1   g567(.A1(G301), .A2(new_n984), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n940), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(G286), .B2(G8), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n995), .B(G8), .C1(new_n535), .C2(new_n537), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(new_n961), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT119), .B(G2084), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n964), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1966), .B1(new_n980), .B2(new_n964), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n999), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n996), .A2(new_n998), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  INV_X1    g585(.A(G1966), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n975), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n964), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1005), .B(new_n1009), .C1(new_n1014), .C2(new_n999), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT51), .B1(new_n999), .B2(KEYINPUT123), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n1007), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT55), .B(G8), .C1(new_n516), .C2(new_n526), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n971), .A2(new_n974), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n858), .A2(new_n1026), .A3(new_n977), .ZN(new_n1027));
  INV_X1    g602(.A(new_n960), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n952), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n964), .A2(new_n970), .A3(new_n957), .A4(new_n955), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1024), .A2(new_n1030), .B1(new_n1031), .B2(new_n804), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1023), .B1(new_n1032), .B2(new_n1010), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n952), .B1(new_n971), .B2(new_n974), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n576), .A2(new_n581), .A3(G1976), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT115), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1036), .A3(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1010), .B1(new_n964), .B2(new_n952), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1036), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT116), .B(G1981), .Z(new_n1044));
  AOI211_X1 g619(.A(new_n1044), .B(new_n592), .C1(new_n588), .C2(G651), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n589), .B2(new_n593), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n513), .A2(G61), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1049), .A2(new_n583), .B1(G73), .B2(G543), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n515), .B1(new_n1050), .B2(new_n586), .ZN(new_n1051));
  OAI21_X1  g626(.A(G1981), .B1(new_n1051), .B2(new_n592), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1044), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n589), .A2(new_n593), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1039), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1038), .A2(new_n1042), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1031), .A2(new_n804), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n963), .A2(new_n1024), .A3(new_n964), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1023), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1033), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n984), .A2(new_n991), .A3(new_n992), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n967), .A2(new_n982), .A3(G301), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(KEYINPUT54), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n994), .A2(new_n1019), .A3(new_n1063), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n953), .A2(new_n955), .A3(new_n957), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n569), .A2(KEYINPUT57), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n563), .B2(new_n568), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT121), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1034), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n964), .A2(KEYINPUT120), .A3(new_n952), .ZN(new_n1087));
  AOI21_X1  g662(.A(G2067), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1348), .B1(new_n963), .B2(new_n964), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n611), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1070), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  AND3_X1   g669(.A1(new_n1086), .A2(new_n1087), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1031), .A2(G1996), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n550), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n550), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT61), .B1(new_n1079), .B2(new_n1092), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NOR4_X1   g678(.A1(new_n1088), .A2(new_n1103), .A3(new_n1089), .A4(new_n611), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1103), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n611), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1083), .A4(new_n1092), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1101), .A2(new_n1105), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1068), .B1(new_n1093), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1038), .A2(new_n1042), .A3(new_n1056), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1038), .A2(new_n1056), .A3(new_n1042), .A4(KEYINPUT117), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1062), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n807), .A2(new_n1040), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT118), .Z(new_n1120));
  OAI21_X1  g695(.A(new_n1054), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1121), .A2(new_n1039), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1061), .B1(new_n1060), .B2(G8), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1010), .B(new_n1023), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1014), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1017), .A2(G286), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1033), .A2(new_n1130), .A3(new_n1057), .A4(new_n1062), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n1112), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1127), .A2(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1092), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n898), .B1(new_n1106), .B2(KEYINPUT60), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1098), .A2(new_n1100), .B1(new_n1143), .B2(new_n1108), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1138), .B(new_n1139), .C1(new_n1145), .C2(new_n1068), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n983), .A3(new_n1063), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1135), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n969), .B1(new_n951), .B2(new_n944), .ZN(new_n1151));
  INV_X1    g726(.A(G1996), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n722), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT112), .Z(new_n1154));
  XNOR2_X1  g729(.A(new_n777), .B(new_n780), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1152), .B2(new_n722), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n792), .A2(new_n796), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n792), .A2(new_n796), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1151), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1986), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n600), .B(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1151), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1150), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT46), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT127), .Z(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1155), .B(new_n722), .C1(new_n1168), .C2(G1996), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1151), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT47), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n778), .A2(new_n780), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1025), .B(new_n969), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1161), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1151), .A2(new_n1162), .A3(new_n600), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1172), .B(new_n1175), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1165), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g755(.A1(new_n466), .A2(G227), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n694), .A2(new_n695), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1183), .B1(new_n655), .B2(new_n658), .ZN(new_n1184));
  AND3_X1   g758(.A1(new_n873), .A2(new_n879), .A3(new_n876), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n879), .B1(new_n873), .B2(new_n876), .ZN(new_n1186));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n936), .B2(new_n937), .ZN(G308));
  OAI221_X1 g762(.A(new_n1184), .B1(new_n1186), .B2(new_n1185), .C1(new_n932), .C2(new_n933), .ZN(G225));
endmodule


