

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n463), .B(KEYINPUT48), .ZN(n541) );
  XOR2_X1 U323 ( .A(n373), .B(n372), .Z(n469) );
  XNOR2_X1 U324 ( .A(n448), .B(n447), .ZN(n496) );
  XOR2_X1 U325 ( .A(G50GAT), .B(G148GAT), .Z(n290) );
  XOR2_X1 U326 ( .A(G106GAT), .B(G78GAT), .Z(n420) );
  XNOR2_X1 U327 ( .A(n310), .B(G162GAT), .ZN(n311) );
  XNOR2_X1 U328 ( .A(n366), .B(n290), .ZN(n367) );
  XNOR2_X1 U329 ( .A(n441), .B(n311), .ZN(n316) );
  XNOR2_X1 U330 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U331 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n470) );
  XOR2_X1 U332 ( .A(KEYINPUT36), .B(n561), .Z(n579) );
  XNOR2_X1 U333 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U334 ( .A(n446), .B(KEYINPUT103), .ZN(n447) );
  XOR2_X1 U335 ( .A(n323), .B(n322), .Z(n561) );
  INV_X1 U336 ( .A(KEYINPUT106), .ZN(n449) );
  XNOR2_X1 U337 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n473) );
  XNOR2_X1 U338 ( .A(n449), .B(G36GAT), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n474), .B(n473), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1329GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n292) );
  XNOR2_X1 U342 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U344 ( .A(n293), .B(G211GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G197GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n370) );
  XOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .Z(n312) );
  XNOR2_X1 U348 ( .A(G176GAT), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n296), .B(G64GAT), .ZN(n416) );
  XOR2_X1 U350 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n298) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n348) );
  XNOR2_X1 U353 ( .A(n416), .B(n348), .ZN(n301) );
  XOR2_X1 U354 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U355 ( .A(n396), .B(KEYINPUT93), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n299), .B(KEYINPUT94), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(n312), .B(n302), .Z(n304) );
  NAND2_X1 U359 ( .A1(G226GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U361 ( .A(n370), .B(n305), .Z(n514) );
  XOR2_X1 U362 ( .A(KEYINPUT65), .B(KEYINPUT77), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT9), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n323) );
  XOR2_X1 U365 ( .A(G43GAT), .B(G50GAT), .Z(n309) );
  XNOR2_X1 U366 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n441) );
  AND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .Z(n423) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(n423), .Z(n314) );
  XNOR2_X1 U371 ( .A(G218GAT), .B(n312), .ZN(n313) );
  XOR2_X1 U372 ( .A(n314), .B(n313), .Z(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U374 ( .A(G29GAT), .B(G134GAT), .Z(n337) );
  XOR2_X1 U375 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n318) );
  XNOR2_X1 U376 ( .A(G92GAT), .B(KEYINPUT66), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n337), .B(n319), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(KEYINPUT2), .B(G162GAT), .Z(n325) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(n326), .ZN(n371) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n327), .B(G148GAT), .ZN(n417) );
  XOR2_X1 U386 ( .A(KEYINPUT4), .B(n417), .Z(n329) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n371), .B(n330), .Z(n344) );
  XOR2_X1 U390 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n332) );
  XNOR2_X1 U391 ( .A(KEYINPUT91), .B(KEYINPUT87), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U393 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n334) );
  XNOR2_X1 U394 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U396 ( .A(n336), .B(n335), .Z(n342) );
  XOR2_X1 U397 ( .A(G113GAT), .B(G1GAT), .Z(n433) );
  XOR2_X1 U398 ( .A(KEYINPUT86), .B(G85GAT), .Z(n339) );
  XOR2_X1 U399 ( .A(KEYINPUT0), .B(G127GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(n347), .B(n337), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n433), .B(n340), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n383) );
  INV_X1 U405 ( .A(n514), .ZN(n464) );
  XOR2_X1 U406 ( .A(G120GAT), .B(G99GAT), .Z(n346) );
  XNOR2_X1 U407 ( .A(G113GAT), .B(G190GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n361) );
  XOR2_X1 U409 ( .A(n348), .B(n347), .Z(n350) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(G134GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U412 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n352) );
  NAND2_X1 U413 ( .A1(G227GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U416 ( .A(G71GAT), .B(G183GAT), .Z(n356) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G176GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n357), .B(KEYINPUT20), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n523) );
  NAND2_X1 U422 ( .A1(n464), .A2(n523), .ZN(n374) );
  XOR2_X1 U423 ( .A(n420), .B(KEYINPUT83), .Z(n363) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U426 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n365) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n373) );
  INV_X1 U430 ( .A(n371), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n374), .A2(n469), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT25), .ZN(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT98), .B(n376), .Z(n380) );
  NOR2_X1 U434 ( .A1(n523), .A2(n469), .ZN(n378) );
  XNOR2_X1 U435 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n565) );
  XOR2_X1 U437 ( .A(KEYINPUT27), .B(n514), .Z(n387) );
  NAND2_X1 U438 ( .A1(n565), .A2(n387), .ZN(n538) );
  XOR2_X1 U439 ( .A(n538), .B(KEYINPUT97), .Z(n379) );
  NAND2_X1 U440 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U441 ( .A1(n383), .A2(n381), .ZN(n382) );
  XNOR2_X1 U442 ( .A(KEYINPUT99), .B(n382), .ZN(n390) );
  XNOR2_X1 U443 ( .A(KEYINPUT92), .B(n383), .ZN(n539) );
  INV_X1 U444 ( .A(n539), .ZN(n385) );
  XNOR2_X1 U445 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n384) );
  XOR2_X1 U446 ( .A(n384), .B(n469), .Z(n520) );
  AND2_X1 U447 ( .A1(n385), .A2(n520), .ZN(n386) );
  NAND2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n525) );
  NOR2_X1 U449 ( .A1(n523), .A2(n525), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT95), .B(n388), .Z(n389) );
  NOR2_X1 U451 ( .A1(n390), .A2(n389), .ZN(n476) );
  NOR2_X1 U452 ( .A1(n579), .A2(n476), .ZN(n409) );
  XOR2_X1 U453 ( .A(G78GAT), .B(KEYINPUT14), .Z(n392) );
  XNOR2_X1 U454 ( .A(G211GAT), .B(G64GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n408) );
  XOR2_X1 U456 ( .A(G57GAT), .B(G155GAT), .Z(n394) );
  XNOR2_X1 U457 ( .A(G1GAT), .B(G127GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U459 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U460 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U462 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U466 ( .A(G15GAT), .B(KEYINPUT71), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(G22GAT), .ZN(n440) );
  XNOR2_X1 U468 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n404), .B(KEYINPUT73), .ZN(n422) );
  XNOR2_X1 U470 ( .A(n440), .B(n422), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n532) );
  INV_X1 U473 ( .A(n532), .ZN(n575) );
  NAND2_X1 U474 ( .A1(n409), .A2(n575), .ZN(n410) );
  XOR2_X1 U475 ( .A(KEYINPUT37), .B(n410), .Z(n511) );
  XOR2_X1 U476 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n412) );
  XNOR2_X1 U477 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n427) );
  XNOR2_X1 U479 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n414) );
  AND2_X1 U480 ( .A1(G230GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U482 ( .A(n415), .B(KEYINPUT76), .Z(n419) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U484 ( .A(n419), .B(n418), .Z(n421) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n571) );
  XOR2_X1 U489 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n429) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(G8GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n445) );
  XOR2_X1 U492 ( .A(G197GAT), .B(G141GAT), .Z(n431) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G36GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U496 ( .A1(G229GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U498 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n437) );
  XNOR2_X1 U499 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U501 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U504 ( .A(n445), .B(n444), .Z(n566) );
  INV_X1 U505 ( .A(n566), .ZN(n552) );
  NAND2_X1 U506 ( .A1(n571), .A2(n552), .ZN(n479) );
  NOR2_X1 U507 ( .A1(n511), .A2(n479), .ZN(n448) );
  XNOR2_X1 U508 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n446) );
  NOR2_X1 U509 ( .A1(n514), .A2(n496), .ZN(n451) );
  INV_X1 U510 ( .A(n523), .ZN(n517) );
  XOR2_X1 U511 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n466) );
  NOR2_X1 U512 ( .A1(n575), .A2(n579), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n452), .B(KEYINPUT45), .ZN(n454) );
  AND2_X1 U514 ( .A1(n571), .A2(n566), .ZN(n453) );
  AND2_X1 U515 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT115), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT41), .B(n571), .Z(n543) );
  NOR2_X1 U519 ( .A1(n566), .A2(n543), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  NOR2_X1 U521 ( .A1(n532), .A2(n457), .ZN(n458) );
  INV_X1 U522 ( .A(n561), .ZN(n550) );
  NAND2_X1 U523 ( .A1(n458), .A2(n550), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n541), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n467), .A2(n539), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT64), .B(n468), .Z(n564) );
  NAND2_X1 U530 ( .A1(n469), .A2(n564), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n517), .A2(n472), .ZN(n560) );
  NAND2_X1 U532 ( .A1(n532), .A2(n560), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n561), .A2(n575), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT16), .ZN(n478) );
  INV_X1 U535 ( .A(n476), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n500) );
  NOR2_X1 U537 ( .A1(n479), .A2(n500), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(n480), .Z(n487) );
  NOR2_X1 U539 ( .A1(n487), .A2(n539), .ZN(n481) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n481), .Z(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(n482), .ZN(G1324GAT) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n514), .A2(n487), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U545 ( .A1(n487), .A2(n517), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n520), .A2(n487), .ZN(n488) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n496), .A2(n539), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n517), .A2(n496), .ZN(n494) );
  XNOR2_X1 U556 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n520), .A2(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n543), .ZN(n557) );
  NAND2_X1 U564 ( .A1(n566), .A2(n557), .ZN(n510) );
  OR2_X1 U565 ( .A1(n500), .A2(n510), .ZN(n507) );
  NOR2_X1 U566 ( .A1(n539), .A2(n507), .ZN(n501) );
  XOR2_X1 U567 ( .A(n501), .B(KEYINPUT42), .Z(n502) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n507), .ZN(n503) );
  XOR2_X1 U570 ( .A(KEYINPUT110), .B(n503), .Z(n504) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n507), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n520), .A2(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  OR2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n539), .A2(n519), .ZN(n512) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U581 ( .A(KEYINPUT112), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n514), .A2(n519), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n517), .A2(n519), .ZN(n518) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n541), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n552), .A2(n535), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U596 ( .A1(n535), .A2(n557), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT117), .Z(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n532), .A2(n535), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U604 ( .A1(n535), .A2(n561), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n549) );
  NOR2_X1 U608 ( .A1(n566), .A2(n549), .ZN(n542) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n549), .A2(n543), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n575), .A2(n549), .ZN(n548) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n560), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n578), .A2(n566), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

