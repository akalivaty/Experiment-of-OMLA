

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770;

  AND2_X1 U377 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U378 ( .A(n562), .B(KEYINPUT115), .ZN(n580) );
  XNOR2_X1 U379 ( .A(n407), .B(n359), .ZN(n525) );
  XNOR2_X1 U380 ( .A(G116), .B(KEYINPUT3), .ZN(n412) );
  NAND2_X1 U381 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X2 U382 ( .A1(n422), .A2(n358), .ZN(n526) );
  INV_X2 U383 ( .A(KEYINPUT65), .ZN(n479) );
  XNOR2_X2 U384 ( .A(n515), .B(n514), .ZN(n747) );
  XNOR2_X2 U385 ( .A(n504), .B(n503), .ZN(n515) );
  NAND2_X2 U386 ( .A1(n425), .A2(n424), .ZN(n627) );
  INV_X1 U387 ( .A(G128), .ZN(n480) );
  XNOR2_X1 U388 ( .A(G119), .B(G128), .ZN(n470) );
  NAND2_X2 U389 ( .A1(n575), .A2(n582), .ZN(n398) );
  XNOR2_X2 U390 ( .A(n526), .B(KEYINPUT39), .ZN(n575) );
  XNOR2_X2 U391 ( .A(n508), .B(n357), .ZN(n669) );
  XNOR2_X2 U392 ( .A(n398), .B(KEYINPUT40), .ZN(n769) );
  XOR2_X2 U393 ( .A(G131), .B(KEYINPUT70), .Z(n529) );
  XNOR2_X2 U394 ( .A(n408), .B(n602), .ZN(n608) );
  XNOR2_X2 U395 ( .A(G478), .B(n356), .ZN(n576) );
  INV_X1 U396 ( .A(KEYINPUT0), .ZN(n417) );
  AND2_X1 U397 ( .A1(n371), .A2(n626), .ZN(n424) );
  OR2_X1 U398 ( .A1(n611), .A2(n767), .ZN(n397) );
  OR2_X1 U399 ( .A1(n611), .A2(KEYINPUT66), .ZN(n626) );
  AND2_X1 U400 ( .A1(n376), .A2(n377), .ZN(n374) );
  XNOR2_X1 U401 ( .A(n394), .B(n609), .ZN(n611) );
  NAND2_X1 U402 ( .A1(n450), .A2(n427), .ZN(n700) );
  NOR2_X1 U403 ( .A1(n571), .A2(n570), .ZN(n432) );
  NAND2_X1 U404 ( .A1(n554), .A2(n577), .ZN(n720) );
  XOR2_X1 U405 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U406 ( .A1(n557), .A2(n666), .ZN(n664) );
  XNOR2_X1 U407 ( .A(n478), .B(n477), .ZN(n557) );
  XNOR2_X1 U408 ( .A(n379), .B(n756), .ZN(n740) );
  INV_X2 U409 ( .A(G953), .ZN(n759) );
  BUF_X1 U410 ( .A(n546), .Z(n355) );
  XNOR2_X1 U411 ( .A(n483), .B(G134), .ZN(n463) );
  XNOR2_X1 U412 ( .A(n433), .B(G146), .ZN(n517) );
  INV_X1 U413 ( .A(G125), .ZN(n433) );
  XNOR2_X1 U414 ( .A(KEYINPUT15), .B(G902), .ZN(n631) );
  XNOR2_X1 U415 ( .A(n745), .B(n448), .ZN(n516) );
  XNOR2_X1 U416 ( .A(n500), .B(KEYINPUT74), .ZN(n448) );
  INV_X1 U417 ( .A(KEYINPUT4), .ZN(n482) );
  XNOR2_X1 U418 ( .A(KEYINPUT72), .B(n560), .ZN(n571) );
  XNOR2_X1 U419 ( .A(n412), .B(G119), .ZN(n504) );
  INV_X1 U420 ( .A(KEYINPUT90), .ZN(n588) );
  AND2_X1 U421 ( .A1(n403), .A2(n404), .ZN(n376) );
  INV_X1 U422 ( .A(G237), .ZN(n509) );
  INV_X1 U423 ( .A(G902), .ZN(n510) );
  NAND2_X1 U424 ( .A1(n413), .A2(n415), .ZN(n372) );
  AND2_X1 U425 ( .A1(n414), .A2(KEYINPUT44), .ZN(n413) );
  NAND2_X1 U426 ( .A1(n611), .A2(KEYINPUT66), .ZN(n415) );
  NOR2_X1 U427 ( .A1(n624), .A2(n623), .ZN(n371) );
  INV_X1 U428 ( .A(KEYINPUT108), .ZN(n370) );
  XOR2_X1 U429 ( .A(KEYINPUT106), .B(G140), .Z(n532) );
  XNOR2_X1 U430 ( .A(G113), .B(G122), .ZN(n531) );
  XNOR2_X1 U431 ( .A(n517), .B(KEYINPUT10), .ZN(n436) );
  XNOR2_X1 U432 ( .A(n530), .B(n438), .ZN(n437) );
  XNOR2_X1 U433 ( .A(n528), .B(G104), .ZN(n438) );
  XNOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n533) );
  XOR2_X1 U435 ( .A(KEYINPUT107), .B(KEYINPUT105), .Z(n534) );
  XNOR2_X1 U436 ( .A(n410), .B(n365), .ZN(n653) );
  XNOR2_X1 U437 ( .A(n430), .B(n429), .ZN(n674) );
  INV_X1 U438 ( .A(KEYINPUT103), .ZN(n429) );
  NOR2_X1 U439 ( .A1(n740), .A2(G902), .ZN(n478) );
  XNOR2_X1 U440 ( .A(n486), .B(n436), .ZN(n756) );
  XNOR2_X1 U441 ( .A(KEYINPUT24), .B(KEYINPUT99), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n516), .B(n447), .ZN(n488) );
  XNOR2_X1 U443 ( .A(n487), .B(n486), .ZN(n447) );
  XNOR2_X1 U444 ( .A(n416), .B(n523), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n747), .B(n516), .ZN(n416) );
  INV_X1 U446 ( .A(KEYINPUT89), .ZN(n651) );
  INV_X1 U447 ( .A(n720), .ZN(n582) );
  NOR2_X1 U448 ( .A1(n653), .A2(n615), .ZN(n389) );
  NOR2_X1 U449 ( .A1(n604), .A2(n459), .ZN(n453) );
  OR2_X1 U450 ( .A1(n453), .A2(KEYINPUT32), .ZN(n451) );
  XNOR2_X1 U451 ( .A(n601), .B(KEYINPUT22), .ZN(n602) );
  XNOR2_X1 U452 ( .A(n539), .B(n434), .ZN(n577) );
  XNOR2_X1 U453 ( .A(n540), .B(n435), .ZN(n434) );
  NAND2_X1 U454 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U455 ( .A1(n717), .A2(n564), .ZN(n568) );
  OR2_X1 U456 ( .A1(KEYINPUT47), .A2(n659), .ZN(n565) );
  INV_X1 U457 ( .A(KEYINPUT86), .ZN(n399) );
  INV_X1 U458 ( .A(n529), .ZN(n483) );
  XNOR2_X1 U459 ( .A(n483), .B(G134), .ZN(n464) );
  INV_X1 U460 ( .A(KEYINPUT109), .ZN(n456) );
  XOR2_X1 U461 ( .A(KEYINPUT69), .B(G101), .Z(n500) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n527) );
  XNOR2_X1 U463 ( .A(n500), .B(n423), .ZN(n501) );
  XNOR2_X1 U464 ( .A(G137), .B(KEYINPUT5), .ZN(n423) );
  INV_X1 U465 ( .A(n766), .ZN(n446) );
  INV_X1 U466 ( .A(KEYINPUT48), .ZN(n418) );
  NAND2_X1 U467 ( .A1(n390), .A2(n631), .ZN(n407) );
  INV_X1 U468 ( .A(G475), .ZN(n435) );
  XNOR2_X1 U469 ( .A(n485), .B(n484), .ZN(n745) );
  XOR2_X1 U470 ( .A(G104), .B(G107), .Z(n485) );
  XNOR2_X1 U471 ( .A(n541), .B(n369), .ZN(n542) );
  XNOR2_X1 U472 ( .A(G134), .B(G122), .ZN(n541) );
  XNOR2_X1 U473 ( .A(n370), .B(KEYINPUT7), .ZN(n369) );
  XNOR2_X1 U474 ( .A(G116), .B(G107), .ZN(n543) );
  NAND2_X1 U475 ( .A1(n480), .A2(KEYINPUT65), .ZN(n386) );
  XNOR2_X1 U476 ( .A(n437), .B(n436), .ZN(n538) );
  XNOR2_X1 U477 ( .A(n401), .B(n616), .ZN(n719) );
  NOR2_X1 U478 ( .A1(n674), .A2(n615), .ZN(n401) );
  INV_X1 U479 ( .A(n621), .ZN(n667) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(G122), .ZN(n513) );
  XNOR2_X1 U481 ( .A(n382), .B(n380), .ZN(n379) );
  XNOR2_X1 U482 ( .A(n472), .B(n381), .ZN(n380) );
  XNOR2_X1 U483 ( .A(n639), .B(KEYINPUT59), .ZN(n640) );
  XNOR2_X1 U484 ( .A(n390), .B(n694), .ZN(n695) );
  XOR2_X1 U485 ( .A(KEYINPUT94), .B(n642), .Z(n729) );
  AND2_X1 U486 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U487 ( .A(n439), .B(KEYINPUT113), .ZN(n766) );
  NAND2_X1 U488 ( .A1(n440), .A2(n553), .ZN(n439) );
  XNOR2_X1 U489 ( .A(n586), .B(n441), .ZN(n440) );
  XNOR2_X1 U490 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n581), .B(KEYINPUT42), .ZN(n768) );
  NAND2_X1 U492 ( .A1(n405), .A2(n663), .ZN(n404) );
  XNOR2_X1 U493 ( .A(n574), .B(n406), .ZN(n405) );
  XNOR2_X1 U494 ( .A(KEYINPUT117), .B(KEYINPUT36), .ZN(n406) );
  NAND2_X1 U495 ( .A1(n388), .A2(n598), .ZN(n387) );
  XNOR2_X1 U496 ( .A(n389), .B(n364), .ZN(n388) );
  NAND2_X1 U497 ( .A1(n454), .A2(n449), .ZN(n427) );
  AND2_X1 U498 ( .A1(n453), .A2(KEYINPUT32), .ZN(n449) );
  NAND2_X1 U499 ( .A1(n580), .A2(n596), .ZN(n717) );
  XNOR2_X1 U500 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U501 ( .A(n669), .B(n366), .ZN(n603) );
  OR2_X1 U502 ( .A1(G902), .A2(n736), .ZN(n356) );
  XNOR2_X1 U503 ( .A(G472), .B(KEYINPUT76), .ZN(n357) );
  XNOR2_X1 U504 ( .A(KEYINPUT38), .B(n553), .ZN(n358) );
  AND2_X1 U505 ( .A1(n524), .A2(G210), .ZN(n359) );
  AND2_X1 U506 ( .A1(n600), .A2(n599), .ZN(n360) );
  INV_X1 U507 ( .A(n570), .ZN(n458) );
  BUF_X1 U508 ( .A(n589), .Z(n663) );
  XOR2_X1 U509 ( .A(G137), .B(G140), .Z(n486) );
  NOR2_X1 U510 ( .A1(n597), .A2(n553), .ZN(n361) );
  AND2_X1 U511 ( .A1(n446), .A2(n587), .ZN(n362) );
  AND2_X1 U512 ( .A1(n446), .A2(n728), .ZN(n363) );
  XNOR2_X1 U513 ( .A(KEYINPUT34), .B(KEYINPUT84), .ZN(n364) );
  XNOR2_X1 U514 ( .A(KEYINPUT33), .B(KEYINPUT75), .ZN(n365) );
  XOR2_X1 U515 ( .A(n569), .B(KEYINPUT6), .Z(n366) );
  XOR2_X1 U516 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n367) );
  AND2_X1 U517 ( .A1(n610), .A2(KEYINPUT92), .ZN(n368) );
  NAND2_X1 U518 ( .A1(n479), .A2(G128), .ZN(n385) );
  XNOR2_X1 U519 ( .A(n507), .B(n488), .ZN(n730) );
  NAND2_X1 U520 ( .A1(n426), .A2(n372), .ZN(n425) );
  XNOR2_X1 U521 ( .A(n373), .B(KEYINPUT71), .ZN(n421) );
  NAND2_X1 U522 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X1 U523 ( .A(n378), .B(n399), .ZN(n375) );
  NAND2_X1 U524 ( .A1(n402), .A2(n568), .ZN(n377) );
  NAND2_X1 U525 ( .A1(n556), .A2(n555), .ZN(n378) );
  NAND2_X1 U526 ( .A1(n547), .A2(G221), .ZN(n382) );
  XNOR2_X2 U527 ( .A(n383), .B(G469), .ZN(n391) );
  OR2_X2 U528 ( .A1(n730), .A2(G902), .ZN(n383) );
  XNOR2_X2 U529 ( .A(n393), .B(G146), .ZN(n507) );
  XNOR2_X2 U530 ( .A(n546), .B(n482), .ZN(n522) );
  XNOR2_X2 U531 ( .A(n384), .B(n481), .ZN(n546) );
  XNOR2_X2 U532 ( .A(n387), .B(KEYINPUT35), .ZN(n767) );
  NAND2_X1 U533 ( .A1(n391), .A2(n664), .ZN(n489) );
  XNOR2_X1 U534 ( .A(n391), .B(KEYINPUT1), .ZN(n589) );
  NAND2_X1 U535 ( .A1(n561), .A2(n391), .ZN(n562) );
  XNOR2_X1 U536 ( .A(n393), .B(n392), .ZN(n761) );
  INV_X1 U537 ( .A(n756), .ZN(n392) );
  NAND2_X2 U538 ( .A1(n462), .A2(n461), .ZN(n393) );
  NAND2_X1 U539 ( .A1(n396), .A2(n714), .ZN(n394) );
  XNOR2_X1 U540 ( .A(n395), .B(n418), .ZN(n444) );
  NAND2_X1 U541 ( .A1(n419), .A2(n421), .ZN(n395) );
  NAND2_X1 U542 ( .A1(n739), .A2(G472), .ZN(n705) );
  AND2_X4 U543 ( .A1(n650), .A2(n638), .ZN(n739) );
  INV_X1 U544 ( .A(n700), .ZN(n396) );
  NAND2_X1 U545 ( .A1(n567), .A2(n566), .ZN(n402) );
  XNOR2_X1 U546 ( .A(n420), .B(n367), .ZN(n419) );
  NAND2_X1 U547 ( .A1(n397), .A2(n368), .ZN(n426) );
  NAND2_X1 U548 ( .A1(n769), .A2(n768), .ZN(n420) );
  NAND2_X1 U549 ( .A1(n400), .A2(n617), .ZN(n457) );
  NAND2_X1 U550 ( .A1(n719), .A2(n710), .ZN(n400) );
  NAND2_X1 U551 ( .A1(n568), .A2(KEYINPUT87), .ZN(n403) );
  INV_X1 U552 ( .A(n404), .ZN(n725) );
  INV_X1 U553 ( .A(n669), .ZN(n570) );
  NOR2_X1 U554 ( .A1(n603), .A2(n571), .ZN(n585) );
  NAND2_X1 U555 ( .A1(n525), .A2(n654), .ZN(n572) );
  NAND2_X1 U556 ( .A1(n431), .A2(n360), .ZN(n408) );
  XNOR2_X2 U557 ( .A(n409), .B(n417), .ZN(n431) );
  NAND2_X2 U558 ( .A1(n596), .A2(n595), .ZN(n409) );
  NAND2_X1 U559 ( .A1(n460), .A2(n459), .ZN(n410) );
  NAND2_X1 U560 ( .A1(n411), .A2(n628), .ZN(n629) );
  NAND2_X1 U561 ( .A1(n411), .A2(n757), .ZN(n646) );
  NAND2_X1 U562 ( .A1(n411), .A2(n759), .ZN(n753) );
  XNOR2_X2 U563 ( .A(n627), .B(KEYINPUT45), .ZN(n411) );
  NAND2_X1 U564 ( .A1(n767), .A2(KEYINPUT92), .ZN(n414) );
  INV_X1 U565 ( .A(n431), .ZN(n615) );
  XNOR2_X2 U566 ( .A(n572), .B(n563), .ZN(n596) );
  NAND2_X1 U567 ( .A1(n422), .A2(n361), .ZN(n701) );
  XNOR2_X2 U568 ( .A(n442), .B(KEYINPUT81), .ZN(n422) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n455) );
  XNOR2_X1 U570 ( .A(n445), .B(n588), .ZN(n628) );
  NAND2_X1 U571 ( .A1(n608), .A2(n455), .ZN(n452) );
  NAND2_X1 U572 ( .A1(n428), .A2(n708), .ZN(n623) );
  XNOR2_X1 U573 ( .A(n457), .B(n456), .ZN(n428) );
  NAND2_X1 U574 ( .A1(n460), .A2(n458), .ZN(n430) );
  NOR2_X1 U575 ( .A1(n512), .A2(n558), .ZN(n443) );
  NAND2_X1 U576 ( .A1(n669), .A2(n654), .ZN(n511) );
  NAND2_X1 U577 ( .A1(n454), .A2(n603), .ZN(n618) );
  XNOR2_X1 U578 ( .A(n432), .B(KEYINPUT28), .ZN(n561) );
  NAND2_X1 U579 ( .A1(n646), .A2(n630), .ZN(n632) );
  AND2_X1 U580 ( .A1(n444), .A2(n363), .ZN(n757) );
  NAND2_X1 U581 ( .A1(n499), .A2(n443), .ZN(n442) );
  NAND2_X1 U582 ( .A1(n444), .A2(n362), .ZN(n445) );
  INV_X1 U583 ( .A(n608), .ZN(n454) );
  INV_X1 U584 ( .A(n603), .ZN(n459) );
  XNOR2_X2 U585 ( .A(n590), .B(KEYINPUT79), .ZN(n460) );
  NAND2_X1 U586 ( .A1(n522), .A2(n463), .ZN(n461) );
  OR2_X2 U587 ( .A1(n522), .A2(n464), .ZN(n462) );
  XNOR2_X1 U588 ( .A(n507), .B(n506), .ZN(n702) );
  BUF_X1 U589 ( .A(n730), .Z(n732) );
  AND2_X1 U590 ( .A1(n685), .A2(n684), .ZN(n465) );
  AND2_X1 U591 ( .A1(n527), .A2(G210), .ZN(n466) );
  XNOR2_X1 U592 ( .A(n501), .B(n466), .ZN(n505) );
  INV_X1 U593 ( .A(KEYINPUT114), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n515), .B(n505), .ZN(n506) );
  INV_X1 U595 ( .A(n525), .ZN(n553) );
  BUF_X1 U596 ( .A(n719), .Z(n723) );
  XNOR2_X1 U597 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n644) );
  NAND2_X1 U598 ( .A1(n631), .A2(G234), .ZN(n467) );
  XNOR2_X1 U599 ( .A(n467), .B(KEYINPUT20), .ZN(n474) );
  AND2_X1 U600 ( .A1(n474), .A2(G221), .ZN(n469) );
  XNOR2_X1 U601 ( .A(KEYINPUT101), .B(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U602 ( .A(n469), .B(n468), .ZN(n666) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(G110), .Z(n471) );
  XNOR2_X1 U604 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U605 ( .A1(G234), .A2(n759), .ZN(n473) );
  XOR2_X1 U606 ( .A(KEYINPUT8), .B(n473), .Z(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT25), .B(KEYINPUT100), .Z(n476) );
  NAND2_X1 U608 ( .A1(G217), .A2(n474), .ZN(n475) );
  XNOR2_X1 U609 ( .A(n476), .B(n475), .ZN(n477) );
  INV_X1 U610 ( .A(G143), .ZN(n481) );
  XNOR2_X1 U611 ( .A(KEYINPUT95), .B(G110), .ZN(n484) );
  NAND2_X1 U612 ( .A1(G227), .A2(n759), .ZN(n487) );
  XNOR2_X2 U613 ( .A(n489), .B(KEYINPUT102), .ZN(n612) );
  XNOR2_X1 U614 ( .A(n612), .B(n490), .ZN(n499) );
  NAND2_X1 U615 ( .A1(G234), .A2(G237), .ZN(n491) );
  XNOR2_X1 U616 ( .A(n491), .B(KEYINPUT14), .ZN(n495) );
  NAND2_X1 U617 ( .A1(G952), .A2(n495), .ZN(n492) );
  XNOR2_X1 U618 ( .A(KEYINPUT96), .B(n492), .ZN(n683) );
  NOR2_X1 U619 ( .A1(G953), .A2(n683), .ZN(n494) );
  INV_X1 U620 ( .A(KEYINPUT97), .ZN(n493) );
  XNOR2_X1 U621 ( .A(n494), .B(n493), .ZN(n594) );
  NAND2_X1 U622 ( .A1(G902), .A2(n495), .ZN(n592) );
  NOR2_X1 U623 ( .A1(G900), .A2(n592), .ZN(n496) );
  NAND2_X1 U624 ( .A1(G953), .A2(n496), .ZN(n497) );
  XNOR2_X1 U625 ( .A(KEYINPUT111), .B(n497), .ZN(n498) );
  NOR2_X1 U626 ( .A1(n594), .A2(n498), .ZN(n558) );
  INV_X1 U627 ( .A(KEYINPUT73), .ZN(n502) );
  XNOR2_X1 U628 ( .A(n502), .B(G113), .ZN(n503) );
  NAND2_X1 U629 ( .A1(n702), .A2(n510), .ZN(n508) );
  NAND2_X1 U630 ( .A1(n510), .A2(n509), .ZN(n524) );
  NAND2_X1 U631 ( .A1(n524), .A2(G214), .ZN(n654) );
  XNOR2_X1 U632 ( .A(KEYINPUT30), .B(n511), .ZN(n512) );
  XNOR2_X1 U633 ( .A(n513), .B(KEYINPUT77), .ZN(n514) );
  XOR2_X1 U634 ( .A(KEYINPUT18), .B(n517), .Z(n520) );
  NAND2_X1 U635 ( .A1(G224), .A2(n759), .ZN(n518) );
  XNOR2_X1 U636 ( .A(n518), .B(KEYINPUT17), .ZN(n519) );
  XNOR2_X1 U637 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U638 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U639 ( .A1(G214), .A2(n527), .ZN(n528) );
  XNOR2_X1 U640 ( .A(G143), .B(n529), .ZN(n530) );
  XNOR2_X1 U641 ( .A(n532), .B(n531), .ZN(n536) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U643 ( .A(n536), .B(n535), .Z(n537) );
  XNOR2_X1 U644 ( .A(n538), .B(n537), .ZN(n639) );
  NOR2_X1 U645 ( .A1(G902), .A2(n639), .ZN(n539) );
  INV_X1 U646 ( .A(KEYINPUT13), .ZN(n540) );
  INV_X1 U647 ( .A(n577), .ZN(n550) );
  XOR2_X1 U648 ( .A(n542), .B(KEYINPUT9), .Z(n544) );
  XNOR2_X1 U649 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U650 ( .A(n355), .B(n545), .Z(n549) );
  NAND2_X1 U651 ( .A1(G217), .A2(n547), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n549), .B(n548), .ZN(n736) );
  NAND2_X1 U653 ( .A1(n550), .A2(n576), .ZN(n722) );
  INV_X1 U654 ( .A(n722), .ZN(n551) );
  NAND2_X1 U655 ( .A1(n575), .A2(n551), .ZN(n728) );
  NAND2_X1 U656 ( .A1(KEYINPUT2), .A2(n728), .ZN(n552) );
  XNOR2_X1 U657 ( .A(KEYINPUT85), .B(n552), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n576), .A2(n577), .ZN(n597) );
  XNOR2_X1 U659 ( .A(n701), .B(KEYINPUT88), .ZN(n556) );
  INV_X1 U660 ( .A(n576), .ZN(n554) );
  NAND2_X1 U661 ( .A1(n722), .A2(n720), .ZN(n617) );
  INV_X1 U662 ( .A(n617), .ZN(n659) );
  NAND2_X1 U663 ( .A1(n659), .A2(KEYINPUT47), .ZN(n555) );
  INV_X1 U664 ( .A(n557), .ZN(n621) );
  NOR2_X1 U665 ( .A1(n558), .A2(n666), .ZN(n559) );
  NAND2_X1 U666 ( .A1(n557), .A2(n559), .ZN(n560) );
  XNOR2_X1 U667 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n563) );
  XNOR2_X1 U668 ( .A(KEYINPUT87), .B(KEYINPUT47), .ZN(n564) );
  XNOR2_X1 U669 ( .A(KEYINPUT78), .B(n565), .ZN(n567) );
  INV_X1 U670 ( .A(n717), .ZN(n566) );
  INV_X1 U671 ( .A(n663), .ZN(n606) );
  INV_X1 U672 ( .A(KEYINPUT110), .ZN(n569) );
  NOR2_X1 U673 ( .A1(n720), .A2(n572), .ZN(n573) );
  NAND2_X1 U674 ( .A1(n585), .A2(n573), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n358), .A2(n654), .ZN(n658) );
  NOR2_X1 U676 ( .A1(n577), .A2(n576), .ZN(n600) );
  INV_X1 U677 ( .A(n600), .ZN(n656) );
  NOR2_X1 U678 ( .A1(n658), .A2(n656), .ZN(n579) );
  XOR2_X1 U679 ( .A(KEYINPUT116), .B(KEYINPUT41), .Z(n578) );
  XNOR2_X1 U680 ( .A(n579), .B(n578), .ZN(n684) );
  NAND2_X1 U681 ( .A1(n684), .A2(n580), .ZN(n581) );
  NAND2_X1 U682 ( .A1(n582), .A2(n654), .ZN(n583) );
  NOR2_X1 U683 ( .A1(n663), .A2(n583), .ZN(n584) );
  NAND2_X1 U684 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U685 ( .A1(n589), .A2(n664), .ZN(n590) );
  NOR2_X1 U686 ( .A1(G898), .A2(n759), .ZN(n591) );
  XOR2_X1 U687 ( .A(KEYINPUT98), .B(n591), .Z(n748) );
  NOR2_X1 U688 ( .A1(n748), .A2(n592), .ZN(n593) );
  OR2_X1 U689 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U690 ( .A(n597), .B(KEYINPUT83), .ZN(n598) );
  INV_X1 U691 ( .A(n666), .ZN(n599) );
  INV_X1 U692 ( .A(KEYINPUT67), .ZN(n601) );
  NAND2_X1 U693 ( .A1(n663), .A2(n667), .ZN(n604) );
  AND2_X1 U694 ( .A1(n570), .A2(n667), .ZN(n605) );
  NAND2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n607) );
  OR2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n714) );
  INV_X1 U697 ( .A(KEYINPUT93), .ZN(n609) );
  INV_X1 U698 ( .A(KEYINPUT66), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n625), .A2(KEYINPUT44), .ZN(n610) );
  NOR2_X1 U700 ( .A1(n767), .A2(KEYINPUT92), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n612), .A2(n458), .ZN(n614) );
  INV_X1 U702 ( .A(n615), .ZN(n613) );
  NAND2_X1 U703 ( .A1(n614), .A2(n613), .ZN(n710) );
  XNOR2_X1 U704 ( .A(KEYINPUT31), .B(KEYINPUT104), .ZN(n616) );
  NOR2_X1 U705 ( .A1(n618), .A2(n663), .ZN(n620) );
  INV_X1 U706 ( .A(KEYINPUT91), .ZN(n619) );
  XNOR2_X1 U707 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n708) );
  XNOR2_X2 U709 ( .A(n629), .B(KEYINPUT80), .ZN(n650) );
  NAND2_X1 U710 ( .A1(KEYINPUT68), .A2(KEYINPUT2), .ZN(n630) );
  INV_X1 U711 ( .A(n631), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n632), .A2(n633), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n633), .A2(KEYINPUT2), .ZN(n635) );
  INV_X1 U714 ( .A(KEYINPUT68), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n739), .A2(G475), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n759), .A2(G952), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n729), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(G60) );
  BUF_X1 U721 ( .A(n646), .Z(n648) );
  INV_X1 U722 ( .A(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(n688) );
  NOR2_X1 U726 ( .A1(n358), .A2(n654), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U728 ( .A(KEYINPUT121), .B(n657), .Z(n661) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U731 ( .A1(n653), .A2(n662), .ZN(n679) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT50), .B(n665), .Z(n672) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT49), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n670), .A2(n458), .ZN(n671) );
  NAND2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n684), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT120), .B(n677), .Z(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U743 ( .A(n680), .B(KEYINPUT52), .ZN(n681) );
  XNOR2_X1 U744 ( .A(KEYINPUT122), .B(n681), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n686) );
  INV_X1 U746 ( .A(n653), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n686), .A2(n465), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n689), .A2(n759), .ZN(n693) );
  XOR2_X1 U749 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n691) );
  INV_X1 U750 ( .A(KEYINPUT124), .ZN(n690) );
  XNOR2_X1 U751 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n693), .B(n692), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n739), .A2(G210), .ZN(n696) );
  XOR2_X1 U754 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n694) );
  XNOR2_X1 U755 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U756 ( .A1(n697), .A2(n729), .ZN(n699) );
  INV_X1 U757 ( .A(KEYINPUT56), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n699), .B(n698), .ZN(G51) );
  XOR2_X1 U759 ( .A(n700), .B(G119), .Z(G21) );
  XNOR2_X1 U760 ( .A(n701), .B(G143), .ZN(G45) );
  XOR2_X1 U761 ( .A(KEYINPUT118), .B(KEYINPUT62), .Z(n703) );
  XNOR2_X1 U762 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U763 ( .A1(n706), .A2(n729), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n707), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U765 ( .A(G101), .B(n708), .ZN(G3) );
  NOR2_X1 U766 ( .A1(n720), .A2(n710), .ZN(n709) );
  XOR2_X1 U767 ( .A(G104), .B(n709), .Z(G6) );
  NOR2_X1 U768 ( .A1(n722), .A2(n710), .ZN(n712) );
  XNOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(G107), .B(n713), .ZN(G9) );
  XNOR2_X1 U772 ( .A(G110), .B(n714), .ZN(G12) );
  NOR2_X1 U773 ( .A1(n717), .A2(n722), .ZN(n716) );
  XNOR2_X1 U774 ( .A(G128), .B(KEYINPUT29), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n716), .B(n715), .ZN(G30) );
  NOR2_X1 U776 ( .A1(n717), .A2(n720), .ZN(n718) );
  XOR2_X1 U777 ( .A(G146), .B(n718), .Z(G48) );
  NOR2_X1 U778 ( .A1(n723), .A2(n720), .ZN(n721) );
  XOR2_X1 U779 ( .A(G113), .B(n721), .Z(G15) );
  NOR2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U781 ( .A(G116), .B(n724), .Z(G18) );
  XOR2_X1 U782 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n727) );
  XNOR2_X1 U783 ( .A(G125), .B(n725), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n727), .B(n726), .ZN(G27) );
  XNOR2_X1 U785 ( .A(G134), .B(n728), .ZN(G36) );
  INV_X1 U786 ( .A(n729), .ZN(n743) );
  NAND2_X1 U787 ( .A1(n739), .A2(G469), .ZN(n734) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n731) );
  XNOR2_X1 U789 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U790 ( .A1(n743), .A2(n735), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n739), .A2(G478), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n736), .B(n737), .ZN(n738) );
  NOR2_X1 U793 ( .A1(n743), .A2(n738), .ZN(G63) );
  NAND2_X1 U794 ( .A1(n739), .A2(G217), .ZN(n742) );
  XNOR2_X1 U795 ( .A(n740), .B(KEYINPUT126), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n742), .B(n741), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(G66) );
  XNOR2_X1 U798 ( .A(G101), .B(n745), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n755) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U805 ( .A(n755), .B(n754), .Z(G69) );
  INV_X1 U806 ( .A(n761), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U809 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U813 ( .A(G140), .B(n766), .Z(G42) );
  XOR2_X1 U814 ( .A(n767), .B(G122), .Z(G24) );
  XNOR2_X1 U815 ( .A(G137), .B(n768), .ZN(G39) );
  BUF_X1 U816 ( .A(n769), .Z(n770) );
  XNOR2_X1 U817 ( .A(G131), .B(n770), .ZN(G33) );
endmodule

