//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n463), .A2(new_n464), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT65), .A4(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(G126), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n462), .A2(KEYINPUT66), .A3(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n462), .A2(KEYINPUT66), .A3(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n492), .B(new_n494), .C1(new_n496), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI211_X1 g078(.A(G50), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G50), .A4(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(new_n508), .B2(new_n509), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT68), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n521), .A2(new_n522), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n508), .B2(new_n509), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n503), .A2(new_n502), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n536), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n533), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n507), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n510), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n545), .A2(new_n546), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n545), .A2(new_n551), .B1(new_n540), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n535), .A2(G43), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(KEYINPUT70), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n507), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n550), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AOI211_X1 g138(.A(KEYINPUT71), .B(new_n561), .C1(new_n555), .C2(new_n558), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT72), .Z(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n535), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n517), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n523), .B2(G91), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  OAI21_X1  g156(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n535), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n530), .A2(new_n510), .A3(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  OAI211_X1 g160(.A(G48), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n540), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G61), .B1(new_n515), .B2(new_n516), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n507), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n507), .B1(new_n596), .B2(KEYINPUT73), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT73), .B2(new_n596), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n545), .A2(new_n599), .B1(new_n540), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n601), .A2(KEYINPUT74), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(KEYINPUT74), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n540), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n609), .A2(KEYINPUT75), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n606), .B1(new_n618), .B2(new_n605), .ZN(G284));
  XOR2_X1   g194(.A(G284), .B(KEYINPUT76), .Z(G321));
  OR3_X1    g195(.A1(G168), .A2(KEYINPUT77), .A3(new_n605), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT77), .B1(G168), .B2(new_n605), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n573), .A2(new_n577), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n621), .B(new_n622), .C1(G868), .C2(new_n623), .ZN(G297));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(G868), .C2(new_n623), .ZN(G280));
  XOR2_X1   g200(.A(KEYINPUT78), .B(G559), .Z(new_n626));
  OAI21_X1  g201(.A(new_n618), .B1(G860), .B2(new_n626), .ZN(G148));
  INV_X1    g202(.A(new_n565), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n605), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n618), .A2(new_n626), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n629), .B1(new_n631), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n493), .A2(new_n469), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n478), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n462), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n493), .A2(new_n462), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n641), .B1(new_n642), .B2(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n639), .A2(new_n640), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(KEYINPUT82), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(KEYINPUT82), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n638), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n647), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n682), .A2(new_n687), .A3(new_n685), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n690));
  AOI211_X1 g265(.A(new_n686), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(new_n693), .ZN(new_n698));
  INV_X1    g273(.A(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n697), .B2(new_n700), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G23), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT86), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT86), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n705), .A2(G6), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n592), .B2(new_n705), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT85), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n711), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT34), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n718), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NOR2_X1   g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n474), .A2(G131), .B1(G119), .B2(new_n478), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G1986), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n705), .A2(G24), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G290), .B2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n738), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n724), .A2(new_n726), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT36), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n727), .A2(G33), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n645), .ZN(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G127), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n473), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(G2105), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n727), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2072), .ZN(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  NOR2_X1   g333(.A1(G164), .A2(new_n727), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G27), .B2(new_n727), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n727), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n474), .A2(G140), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n462), .A2(G116), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n478), .A2(KEYINPUT88), .A3(G128), .ZN(new_n767));
  AOI21_X1  g342(.A(KEYINPUT88), .B1(new_n478), .B2(G128), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n764), .B1(new_n765), .B2(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n763), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT89), .B(G2067), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT30), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G160), .A2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n778), .B1(new_n727), .B2(new_n646), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n705), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n705), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n785), .B1(G1961), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n761), .A2(new_n772), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(G29), .A2(G32), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n469), .A2(G105), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n478), .A2(G129), .ZN(new_n796));
  INV_X1    g371(.A(G141), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n645), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n790), .B1(new_n800), .B2(new_n727), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT27), .B(G1996), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n801), .A2(KEYINPUT92), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n789), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n705), .A2(G20), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT23), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G1956), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n810), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G1956), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2090), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n727), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n727), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT29), .Z(new_n820));
  OAI211_X1 g395(.A(new_n812), .B(new_n816), .C1(new_n817), .C2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(G4), .A2(G16), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n618), .B2(G16), .ZN(new_n826));
  INV_X1    g401(.A(G1348), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n807), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n787), .A2(G1961), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n784), .B2(new_n783), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n801), .B2(new_n802), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT93), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n705), .A2(G19), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT87), .Z(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n628), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1341), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n838), .A3(new_n817), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n760), .A2(new_n758), .ZN(new_n840));
  INV_X1    g415(.A(G1966), .ZN(new_n841));
  NOR2_X1   g416(.A1(G168), .A2(new_n705), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n705), .B2(G21), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n841), .B2(new_n843), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n838), .B1(new_n820), .B2(new_n817), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n833), .A2(new_n837), .A3(new_n839), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n829), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n745), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n745), .B2(new_n849), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(G311));
  NAND2_X1  g428(.A1(new_n745), .A2(new_n849), .ZN(G150));
  AOI22_X1  g429(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n507), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n545), .A2(new_n857), .B1(new_n540), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n563), .B2(new_n564), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n559), .A2(new_n562), .A3(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n618), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n861), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  INV_X1    g448(.A(new_n799), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(new_n755), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n800), .B2(new_n755), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n500), .A2(KEYINPUT99), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n487), .A2(new_n491), .B1(new_n478), .B2(G126), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT4), .B1(new_n473), .B2(new_n495), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n493), .A2(new_n497), .A3(new_n498), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n769), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n876), .A2(new_n885), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n735), .A2(new_n635), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n735), .A2(new_n635), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n474), .A2(G142), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT100), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  INV_X1    g468(.A(G118), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(G2105), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G130), .B2(new_n478), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n890), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n886), .A2(new_n887), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n898), .B(KEYINPUT101), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n886), .A2(new_n887), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n482), .B(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT98), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n646), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  INV_X1    g485(.A(new_n904), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n902), .A2(new_n903), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n909), .A2(new_n910), .A3(new_n913), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  NAND2_X1  g494(.A1(G303), .A2(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(G166), .A2(new_n707), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(new_n592), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G290), .B(G305), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n920), .A3(new_n921), .ZN(new_n926));
  XOR2_X1   g501(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n927));
  AND3_X1   g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n924), .A2(new_n926), .B1(new_n929), .B2(KEYINPUT42), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n623), .A2(new_n609), .A3(new_n613), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n614), .A2(G299), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT104), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n614), .A2(G299), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n609), .A2(new_n613), .B1(new_n573), .B2(new_n577), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT41), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n935), .A3(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n553), .A2(new_n554), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT70), .B1(new_n556), .B2(new_n557), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n562), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT71), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n559), .A2(new_n550), .A3(new_n562), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n860), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n863), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n630), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n631), .A2(new_n864), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n941), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n937), .A2(new_n938), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n931), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n936), .A2(new_n940), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n950), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n954), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT106), .B1(new_n962), .B2(new_n931), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n928), .A2(new_n930), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n954), .A4(new_n961), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(KEYINPUT107), .A3(new_n931), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n958), .A2(new_n963), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G868), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT108), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n861), .A2(new_n605), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(new_n972), .A3(G868), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(G295));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(G331));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n924), .A2(new_n926), .ZN(new_n977));
  XNOR2_X1  g552(.A(G168), .B(G171), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n947), .B2(new_n948), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n953), .ZN(new_n980));
  XNOR2_X1  g555(.A(G168), .B(G301), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n862), .A2(new_n981), .A3(new_n863), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n862), .A2(new_n981), .A3(KEYINPUT109), .A4(new_n863), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n979), .A2(new_n982), .B1(new_n935), .B2(new_n939), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n977), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n977), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n979), .A2(new_n982), .A3(new_n953), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n984), .A2(new_n985), .B1(new_n864), .B2(new_n978), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(new_n941), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n992), .A3(new_n910), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n988), .A2(new_n992), .A3(new_n995), .A4(new_n910), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n976), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n992), .A2(new_n910), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n991), .B2(new_n941), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n977), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT43), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT44), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n976), .B1(new_n998), .B2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(G397));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n1008));
  OAI21_X1  g583(.A(G1981), .B1(new_n588), .B2(new_n591), .ZN(new_n1009));
  INV_X1    g584(.A(G61), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n521), .B2(new_n522), .ZN(new_n1011));
  INV_X1    g586(.A(new_n590), .ZN(new_n1012));
  OAI21_X1  g587(.A(G651), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n530), .A2(new_n510), .A3(G86), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n586), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1009), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT49), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n878), .B2(new_n881), .ZN(new_n1021));
  INV_X1    g596(.A(G40), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n467), .A2(new_n471), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n500), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n707), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1019), .A2(new_n1024), .B1(KEYINPUT52), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1026), .A2(G8), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT114), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1024), .A2(new_n1034), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G160), .A2(G40), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n496), .A2(new_n499), .ZN(new_n1039));
  INV_X1    g614(.A(new_n486), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT65), .B1(new_n1040), .B2(new_n490), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n485), .A2(new_n486), .A3(new_n484), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n494), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1025), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(G1384), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n877), .A2(new_n883), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1023), .B1(new_n1021), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT50), .B(G1384), .C1(new_n878), .C2(new_n881), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n817), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1020), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n527), .A2(G8), .A3(new_n528), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n527), .A2(KEYINPUT55), .A3(G8), .A4(new_n528), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1037), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1021), .A2(new_n1051), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1023), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G2090), .B1(new_n1066), .B2(KEYINPUT116), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .A4(new_n1023), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1049), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1063), .B1(new_n1070), .B2(new_n1020), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n500), .A2(new_n1047), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(new_n1023), .C1(new_n1021), .C2(KEYINPUT45), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n841), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1064), .A2(new_n1065), .A3(new_n784), .A4(new_n1023), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G168), .A2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1062), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1037), .A2(KEYINPUT115), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1029), .A2(new_n1036), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1052), .A2(new_n1053), .A3(G2090), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n1049), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1063), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1061), .B(G8), .C1(new_n1049), .C2(new_n1085), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1089), .B(new_n1077), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1079), .A2(new_n1080), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1030), .A3(new_n707), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(G1981), .B2(G305), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1024), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1008), .B1(new_n1092), .B2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT116), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n817), .A3(new_n1069), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1020), .B1(new_n1103), .B2(new_n1050), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(new_n1088), .C1(new_n1104), .C2(new_n1061), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1078), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1080), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1091), .A2(new_n1084), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1100), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  INV_X1    g689(.A(G1961), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1023), .A3(new_n1072), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1046), .A2(new_n1048), .A3(new_n758), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1121), .A2(KEYINPUT122), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1116), .A2(new_n1124), .A3(new_n1120), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1122), .A2(new_n1118), .B1(new_n1066), .B2(new_n1115), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n882), .B1(new_n878), .B2(new_n881), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT45), .B1(new_n1130), .B2(new_n1025), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1023), .A2(new_n1119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1048), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1045), .B1(new_n884), .B2(G1384), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1048), .A4(new_n1132), .ZN(new_n1137));
  AND4_X1   g712(.A1(G301), .A2(new_n1127), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1114), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1062), .A2(new_n1071), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1076), .A2(G168), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1074), .A2(new_n1075), .A3(G168), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G8), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT51), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1144), .A2(KEYINPUT51), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1113), .A2(new_n1139), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1127), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT126), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1127), .A2(new_n1134), .A3(new_n1151), .A4(new_n1137), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(G171), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1123), .A2(G301), .A3(new_n1125), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT125), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1123), .A2(new_n1156), .A3(G301), .A4(new_n1125), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1153), .A2(new_n1155), .A3(KEYINPUT54), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1066), .A2(new_n815), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G299), .B(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1046), .A2(new_n1048), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1054), .A2(G1348), .B1(G2067), .B2(new_n1026), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n618), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G299), .B(KEYINPUT57), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1046), .A2(new_n1048), .A3(new_n1164), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1038), .B1(new_n1044), .B2(KEYINPUT50), .ZN(new_n1171));
  AOI21_X1  g746(.A(G1956), .B1(new_n1171), .B2(new_n1065), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n1173), .B2(new_n1166), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(KEYINPUT121), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1177), .B(KEYINPUT61), .C1(new_n1173), .C2(new_n1166), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n618), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1026), .A2(G2067), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n1066), .B2(new_n827), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n618), .A3(KEYINPUT60), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(G1996), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1046), .A2(new_n1048), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT58), .B(G1341), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1026), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(KEYINPUT119), .A3(new_n565), .ZN(new_n1193));
  XOR2_X1   g768(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1194));
  OR2_X1    g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1173), .A2(new_n1166), .A3(KEYINPUT61), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1187), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1174), .B1(new_n1179), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(G301), .B1(new_n1149), .B2(KEYINPUT126), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1114), .B1(new_n1200), .B2(new_n1152), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1201), .A2(KEYINPUT127), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1148), .A2(new_n1160), .A3(new_n1199), .A4(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1113), .A2(new_n1141), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1147), .A2(KEYINPUT62), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1147), .A2(KEYINPUT62), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1126), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1112), .A2(new_n1203), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1131), .A2(new_n1023), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT111), .Z(new_n1210));
  XOR2_X1   g785(.A(new_n769), .B(G2067), .Z(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT112), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n874), .A2(G1996), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1213), .B1(new_n800), .B2(G1996), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n735), .B(new_n737), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OR2_X1    g792(.A1(G290), .A2(G1986), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(G290), .A2(G1986), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1210), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1222), .B(KEYINPUT113), .Z(new_n1223));
  NAND2_X1  g798(.A1(new_n1208), .A2(new_n1223), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1210), .A2(new_n1219), .ZN(new_n1225));
  OR2_X1    g800(.A1(new_n1225), .A2(KEYINPUT48), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(KEYINPUT48), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1226), .A2(new_n1217), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n735), .A2(new_n737), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1215), .A2(new_n1229), .B1(G2067), .B2(new_n769), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1210), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1210), .A2(new_n1188), .ZN(new_n1233));
  XNOR2_X1  g808(.A(new_n1233), .B(KEYINPUT46), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1210), .B1(new_n874), .B2(new_n1212), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(KEYINPUT47), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT47), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1234), .A2(new_n1238), .A3(new_n1235), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1232), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1224), .A2(new_n1240), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g816(.A1(G227), .A2(new_n460), .ZN(new_n1243));
  OAI21_X1  g817(.A(new_n1243), .B1(new_n702), .B2(new_n703), .ZN(new_n1244));
  NOR2_X1   g818(.A1(new_n1244), .A2(G401), .ZN(new_n1245));
  OAI211_X1 g819(.A(new_n914), .B(new_n1245), .C1(new_n1004), .C2(new_n1005), .ZN(G225));
  INV_X1    g820(.A(G225), .ZN(G308));
endmodule


