//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n204), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n210), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n218), .A2(new_n229), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n213), .A2(new_n214), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n204), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n249), .A2(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G50), .A2(G58), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n204), .B1(new_n255), .B2(new_n222), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n248), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n213), .A2(new_n258), .A3(new_n214), .A4(new_n247), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n257), .B(new_n262), .C1(G50), .C2(new_n258), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G222), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(G1698), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n269), .B1(new_n270), .B2(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n213), .A2(new_n214), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(G274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n281), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(G226), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n263), .B1(new_n288), .B2(G169), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(G179), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n288), .A2(new_n292), .B1(new_n293), .B2(new_n263), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n263), .A2(new_n293), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n287), .B2(new_n296), .ZN(new_n297));
  OR3_X1    g0097(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT10), .B1(new_n294), .B2(new_n297), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n291), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(G226), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n277), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n283), .B1(G238), .B2(new_n285), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n301), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(G190), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n310), .ZN(new_n312));
  OAI21_X1  g0112(.A(G200), .B1(new_n312), .B2(new_n308), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n253), .A2(new_n220), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n250), .A2(new_n270), .B1(new_n204), .B2(G68), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n248), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT68), .ZN(new_n318));
  AOI211_X1 g0118(.A(G68), .B(new_n258), .C1(new_n318), .C2(KEYINPUT12), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(KEYINPUT12), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n317), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n311), .A2(new_n313), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n311), .A2(new_n313), .A3(new_n327), .A4(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(G169), .C1(new_n312), .C2(new_n308), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n309), .A2(new_n310), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(G169), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n250), .B1(new_n204), .B2(new_n270), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n249), .A2(new_n253), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n248), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n261), .A2(G77), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n259), .A2(new_n344), .B1(G77), .B2(new_n258), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n268), .A2(G232), .B1(new_n350), .B2(G107), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n223), .B2(new_n273), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n277), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n283), .B1(G244), .B2(new_n285), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n347), .B(KEYINPUT67), .C1(G169), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT67), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n345), .B1(new_n341), .B2(new_n342), .ZN(new_n358));
  AOI21_X1  g0158(.A(G169), .B1(new_n353), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n332), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(G190), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n358), .C1(new_n292), .C2(new_n355), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n300), .A2(new_n329), .A3(new_n336), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n249), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n261), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n368), .A2(new_n259), .B1(new_n258), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(new_n248), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT70), .B1(new_n348), .B2(new_n349), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n266), .A2(new_n372), .A3(new_n267), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n373), .A3(new_n204), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR4_X1   g0176(.A1(new_n348), .A2(new_n349), .A3(new_n375), .A4(G20), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT71), .A3(G68), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n374), .B2(new_n375), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n222), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G58), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n222), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n370), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n350), .B2(new_n204), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n392), .B2(new_n377), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n369), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n285), .A2(G232), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n282), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n275), .A2(new_n276), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n221), .A2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n271), .B(new_n400), .C1(G223), .C2(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G169), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n398), .A2(new_n403), .A3(new_n332), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT18), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT71), .B1(new_n379), .B2(G68), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n382), .A2(new_n381), .A3(new_n222), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n390), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n395), .A3(new_n248), .ZN(new_n413));
  INV_X1    g0213(.A(new_n369), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(new_n296), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G200), .B2(new_n404), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(new_n408), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n394), .B(new_n370), .C1(new_n384), .C2(new_n390), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(new_n369), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n416), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n409), .A2(new_n419), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n366), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(G20), .B1(G33), .B2(G283), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n265), .A2(G97), .ZN(new_n428));
  INV_X1    g0228(.A(G116), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n427), .A2(new_n428), .B1(G20), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n248), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT20), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n248), .A3(KEYINPUT20), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT82), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n258), .A2(new_n429), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n265), .A2(G1), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n259), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n431), .A2(new_n440), .A3(new_n432), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n443));
  INV_X1    g0243(.A(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(G257), .B(new_n444), .C1(new_n348), .C2(new_n349), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT81), .B(G303), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n443), .B(new_n445), .C1(new_n271), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n277), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G41), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n450), .A2(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G270), .A3(new_n281), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n281), .A2(G274), .A3(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n451), .A2(new_n453), .B1(new_n450), .B2(G41), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n448), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G169), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT83), .B1(new_n442), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(G169), .A4(new_n464), .ZN(new_n469));
  XOR2_X1   g0269(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n470));
  NAND3_X1  g0270(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n464), .A2(G200), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n442), .A2(new_n472), .A3(KEYINPUT85), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n447), .A2(new_n277), .B1(new_n461), .B2(new_n462), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n292), .B1(new_n475), .B2(new_n459), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n476), .B2(new_n467), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(G190), .A3(new_n459), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n464), .A2(KEYINPUT21), .A3(G169), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n448), .A2(G179), .A3(new_n459), .A4(new_n463), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n467), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n471), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n284), .B1(new_n462), .B2(new_n456), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(G257), .B1(new_n462), .B2(new_n461), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n266), .B2(new_n267), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g0289(.A(G1698), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT4), .A2(G244), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n444), .B(new_n492), .C1(new_n348), .C2(new_n349), .ZN(new_n493));
  INV_X1    g0293(.A(G244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n489), .B1(new_n350), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT75), .B1(new_n496), .B2(new_n277), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n266), .B2(new_n267), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n493), .B(new_n491), .C1(new_n498), .C2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n348), .B2(new_n349), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n444), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT75), .B(new_n277), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n486), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT77), .B1(new_n504), .B2(G179), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n485), .A2(G257), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n463), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n277), .B1(new_n499), .B2(new_n501), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT75), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n502), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT77), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n332), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  AND2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g0319(.A1(KEYINPUT6), .A2(G97), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(G107), .ZN(new_n521));
  INV_X1    g0321(.A(G107), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(KEYINPUT73), .A3(KEYINPUT6), .A4(G97), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n518), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT72), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n253), .B2(new_n270), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n252), .A2(KEYINPUT72), .A3(G77), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n524), .A2(G20), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT74), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G107), .B1(new_n392), .B2(new_n377), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n248), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n258), .A2(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n438), .B2(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n486), .A2(new_n508), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n533), .A2(new_n535), .B1(new_n405), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n504), .A2(G200), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n486), .A2(G190), .A3(new_n508), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n514), .A2(new_n537), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n444), .C1(new_n348), .C2(new_n349), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G294), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n277), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n458), .A2(G264), .A3(new_n281), .ZN(new_n547));
  AND4_X1   g0347(.A1(G179), .A2(new_n546), .A3(new_n547), .A4(new_n463), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n485), .A2(G264), .B1(new_n545), .B2(new_n277), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n405), .B1(new_n549), .B2(new_n463), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n547), .A3(new_n463), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G169), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT86), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n204), .B(G87), .C1(new_n348), .C2(new_n349), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n271), .A2(new_n558), .A3(new_n204), .A4(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G116), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n204), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n522), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n560), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n561), .B1(new_n560), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n248), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n258), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n522), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT25), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(G107), .B2(new_n438), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n552), .A2(new_n555), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n438), .A2(G87), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n204), .B1(new_n304), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n517), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n204), .B(G68), .C1(new_n348), .C2(new_n349), .ZN(new_n582));
  INV_X1    g0382(.A(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n577), .B1(new_n250), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n248), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n337), .A2(new_n571), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n576), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n460), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n281), .A2(KEYINPUT78), .A3(G274), .A4(new_n456), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n456), .A2(new_n487), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n590), .A2(new_n591), .B1(new_n281), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n594));
  OAI211_X1 g0394(.A(G238), .B(new_n444), .C1(new_n348), .C2(new_n349), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n562), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n277), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(G190), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n281), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n588), .B(new_n598), .C1(new_n601), .C2(new_n292), .ZN(new_n602));
  INV_X1    g0402(.A(new_n337), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n438), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n586), .A3(new_n587), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT80), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(new_n586), .A3(new_n607), .A4(new_n587), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT79), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n593), .A2(new_n609), .A3(new_n332), .A4(new_n597), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n593), .A2(new_n332), .A3(new_n597), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n593), .A2(new_n597), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n405), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n602), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n549), .A2(G190), .A3(new_n463), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n553), .A2(G200), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n570), .A2(new_n574), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n575), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n426), .A2(new_n484), .A3(new_n541), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(KEYINPUT90), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n362), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n356), .A2(KEYINPUT90), .A3(new_n360), .A4(new_n361), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n329), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n336), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n419), .A2(new_n424), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT89), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n413), .A2(new_n414), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n420), .B1(new_n631), .B2(new_n421), .ZN(new_n632));
  AOI211_X1 g0432(.A(KEYINPUT18), .B(new_n408), .C1(new_n413), .C2(new_n414), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n409), .A2(KEYINPUT89), .A3(new_n423), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n298), .A2(new_n299), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n291), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n504), .A2(KEYINPUT77), .A3(G179), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n512), .B1(new_n511), .B2(new_n332), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n537), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n540), .A2(new_n538), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n612), .B(new_n605), .C1(new_n601), .C2(G169), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n602), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n620), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT87), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n541), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n471), .A2(new_n483), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n575), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n602), .A2(new_n644), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n655), .B(new_n537), .C1(new_n640), .C2(new_n641), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT88), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(KEYINPUT88), .A3(new_n657), .ZN(new_n659));
  INV_X1    g0459(.A(new_n617), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(new_n514), .A3(KEYINPUT26), .A4(new_n537), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n654), .B(new_n644), .C1(new_n658), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n426), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n639), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(G213), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT91), .Z(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT92), .B(G343), .Z(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n442), .ZN(new_n675));
  MUX2_X1   g0475(.A(new_n484), .B(new_n651), .S(new_n675), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n570), .A2(new_n574), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n673), .A2(KEYINPUT93), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT93), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  OR4_X1    g0481(.A1(new_n575), .A2(new_n680), .A3(new_n681), .A4(new_n620), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n575), .A2(new_n673), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n651), .A2(new_n674), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n682), .B2(new_n684), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n575), .A2(new_n674), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n207), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n580), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n216), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n644), .B1(new_n662), .B2(new_n658), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n699), .B(new_n674), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n644), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n656), .B2(KEYINPUT26), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n660), .A2(new_n514), .A3(new_n657), .A4(new_n537), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n705), .C1(new_n647), .C2(new_n652), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n674), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n593), .A2(new_n597), .A3(new_n547), .A4(new_n546), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n536), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT30), .B1(new_n712), .B2(new_n482), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n464), .A2(new_n614), .A3(new_n553), .A4(new_n332), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n511), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n601), .A2(new_n486), .A3(new_n508), .A4(new_n549), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n481), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n464), .A2(new_n614), .A3(new_n332), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n504), .A2(new_n720), .A3(new_n553), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT95), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n718), .A2(new_n717), .A3(new_n481), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n674), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n536), .A2(new_n711), .A3(new_n481), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .B1(new_n511), .B2(new_n714), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n673), .B1(new_n729), .B2(new_n723), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n725), .A2(new_n727), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n541), .A2(new_n621), .A3(new_n484), .A4(new_n674), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT96), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n736), .A3(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n709), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n698), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(G13), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n203), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n693), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n678), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n676), .ZN(new_n747));
  INV_X1    g0547(.A(new_n745), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n275), .B1(new_n204), .B2(G169), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT97), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n204), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n752), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G329), .A2(new_n754), .B1(new_n758), .B2(G311), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n755), .A2(new_n292), .A3(G190), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n761), .A2(G303), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n755), .A2(new_n296), .A3(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n271), .B1(G322), .B2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n759), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n204), .A2(new_n292), .A3(G179), .A4(G190), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n769), .A2(G326), .B1(new_n770), .B2(G283), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n296), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n204), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n767), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n754), .A2(G159), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  INV_X1    g0577(.A(new_n765), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n271), .B1(new_n757), .B2(new_n270), .C1(new_n778), .C2(new_n385), .ZN(new_n779));
  INV_X1    g0579(.A(new_n762), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n222), .B1(new_n768), .B2(new_n220), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n770), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n783), .A2(new_n522), .B1(new_n774), .B2(new_n583), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n760), .A2(new_n579), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n775), .A2(KEYINPUT99), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n750), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n750), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT98), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n692), .A2(new_n350), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G355), .B1(new_n429), .B2(new_n692), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n371), .A2(new_n373), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n692), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n216), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n245), .A2(new_n455), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n748), .B(new_n789), .C1(new_n796), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n676), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n747), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n365), .A2(new_n674), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n659), .A2(new_n661), .ZN(new_n810));
  INV_X1    g0610(.A(new_n658), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n703), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n809), .B1(new_n812), .B2(new_n654), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n673), .B1(new_n812), .B2(new_n654), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n673), .A2(new_n347), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n365), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n624), .A2(new_n625), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n816), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n814), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n738), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n823), .A2(new_n748), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n758), .A2(G159), .B1(G143), .B2(new_n765), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n768), .C1(new_n251), .C2(new_n780), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(new_n799), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G132), .B2(new_n754), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n761), .A2(G50), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n783), .A2(new_n222), .ZN(new_n834));
  INV_X1    g0634(.A(new_n774), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(G58), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n830), .A2(new_n832), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n753), .A2(new_n838), .B1(new_n757), .B2(new_n429), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n271), .B(new_n839), .C1(G294), .C2(new_n765), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n761), .A2(G107), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n769), .A2(G303), .B1(new_n770), .B2(G87), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n835), .A2(G97), .B1(G283), .B2(new_n762), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n750), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n750), .A2(new_n792), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT100), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n748), .B(new_n845), .C1(new_n270), .C2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n819), .B2(new_n792), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n826), .A2(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n742), .A2(new_n203), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n636), .A2(new_n670), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n389), .B1(new_n410), .B2(new_n411), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT16), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n369), .B1(new_n856), .B2(new_n391), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n417), .B1(new_n857), .B2(new_n408), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n671), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n631), .A2(new_n421), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n631), .A2(new_n670), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n417), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n425), .A2(new_n859), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT103), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI211_X1 g0670(.A(KEYINPUT103), .B(KEYINPUT38), .C1(new_n865), .C2(new_n866), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n362), .A2(new_n673), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT102), .Z(new_n874));
  INV_X1    g0674(.A(new_n809), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n663), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n673), .A2(new_n323), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n329), .A2(new_n336), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n329), .B2(new_n336), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n853), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n870), .B2(new_n871), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n862), .B1(new_n636), .B2(new_n628), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n861), .A2(new_n862), .A3(new_n417), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n863), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n867), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n336), .A2(new_n673), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n883), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n709), .A2(new_n426), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n639), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(G330), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n865), .A2(new_n866), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n885), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n902));
  INV_X1    g0702(.A(new_n871), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n730), .B(KEYINPUT31), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n732), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n880), .A2(new_n819), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  AND4_X1   g0708(.A1(KEYINPUT40), .A2(new_n880), .A3(new_n819), .A4(new_n905), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(new_n908), .B1(new_n890), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n426), .A2(new_n905), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n852), .B1(new_n898), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n898), .B2(new_n913), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n916), .A2(G116), .A3(new_n215), .A4(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n386), .A2(new_n216), .A3(new_n270), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n222), .A2(G50), .ZN(new_n921));
  OAI211_X1 g0721(.A(G1), .B(new_n741), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(G367));
  NOR2_X1   g0723(.A1(new_n760), .A2(new_n385), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n774), .A2(new_n222), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(G159), .C2(new_n762), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n753), .A2(new_n828), .B1(new_n757), .B2(new_n220), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n350), .B(new_n927), .C1(G150), .C2(new_n765), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n770), .A2(G77), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n769), .A2(G143), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n760), .A2(new_n429), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT46), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n780), .A2(new_n772), .B1(new_n768), .B2(new_n838), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G97), .B2(new_n770), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n754), .A2(G317), .ZN(new_n936));
  INV_X1    g0736(.A(new_n446), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n758), .A2(G283), .B1(new_n937), .B2(new_n765), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n799), .B1(new_n835), .B2(G107), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n935), .A2(new_n936), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n931), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT105), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n750), .B1(new_n942), .B2(KEYINPUT47), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT47), .B2(new_n942), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n800), .A2(new_n238), .B1(new_n692), .B2(new_n603), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n748), .B1(new_n794), .B2(new_n945), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n674), .A2(new_n588), .A3(new_n644), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n655), .B1(new_n674), .B2(new_n588), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n946), .C1(new_n805), .C2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n533), .A2(new_n535), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n541), .B1(new_n951), .B2(new_n674), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n514), .A2(new_n537), .A3(new_n673), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n690), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n688), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n689), .A2(new_n690), .A3(new_n954), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n690), .A4(new_n954), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n686), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n964), .A3(new_n686), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n687), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT104), .B1(new_n685), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n678), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n677), .B(KEYINPUT104), .C1(new_n685), .C2(new_n970), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n972), .A2(new_n688), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n688), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n739), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n693), .B(KEYINPUT41), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n744), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n949), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT43), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n688), .A2(new_n954), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n643), .A2(new_n575), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n673), .B1(new_n986), .B2(new_n642), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(KEYINPUT42), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n983), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n985), .A2(new_n988), .A3(new_n982), .A4(new_n981), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n686), .A2(new_n955), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n993), .B1(new_n990), .B2(new_n991), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n950), .B1(new_n980), .B2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n695), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n797), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(G107), .B2(new_n207), .ZN(new_n1002));
  AOI211_X1 g0802(.A(G45), .B(new_n1000), .C1(G68), .C2(G77), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n249), .A2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n692), .B(new_n799), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n235), .A2(G45), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n745), .B1(new_n795), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n778), .A2(new_n220), .B1(new_n757), .B2(new_n222), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G150), .B2(new_n754), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n831), .B1(G97), .B2(new_n770), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n835), .A2(new_n603), .B1(new_n769), .B2(G159), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n761), .A2(G77), .B1(new_n367), .B2(new_n762), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n799), .B1(G326), .B2(new_n754), .ZN(new_n1016));
  INV_X1    g0816(.A(G283), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n774), .A2(new_n1017), .B1(new_n760), .B2(new_n772), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n758), .A2(new_n937), .B1(G317), .B2(new_n765), .ZN(new_n1019));
  INV_X1    g0819(.A(G322), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n838), .B2(new_n780), .C1(new_n1020), .C2(new_n768), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1016), .B1(new_n429), .B2(new_n783), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1015), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1009), .B1(new_n1028), .B2(new_n790), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n685), .B2(new_n805), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT106), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n976), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n744), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n976), .A2(new_n738), .A3(new_n709), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n693), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1032), .A2(new_n739), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  AOI22_X1  g0838(.A1(new_n800), .A2(new_n242), .B1(G97), .B2(new_n692), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n748), .B1(new_n794), .B2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n350), .B1(new_n1020), .B2(new_n753), .C1(new_n783), .C2(new_n522), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G283), .B2(new_n761), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT107), .Z(new_n1043));
  OAI22_X1  g0843(.A1(new_n774), .A2(new_n429), .B1(new_n757), .B2(new_n772), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n769), .A2(G317), .B1(G311), .B2(new_n765), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1044), .B(new_n1046), .C1(new_n937), .C2(new_n762), .ZN(new_n1047));
  INV_X1    g0847(.A(G159), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n778), .A2(new_n1048), .B1(new_n768), .B2(new_n251), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n754), .A2(G143), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n799), .C1(new_n249), .C2(new_n757), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n783), .A2(new_n579), .B1(new_n220), .B2(new_n780), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n760), .A2(new_n222), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n774), .A2(new_n270), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1043), .A2(new_n1047), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1040), .B1(new_n750), .B2(new_n1057), .C1(new_n954), .C2(new_n805), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n969), .B2(new_n743), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n968), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n686), .B1(new_n959), .B2(new_n964), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n694), .B1(new_n1062), .B2(new_n1034), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1035), .A2(new_n969), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(G390));
  OAI21_X1  g0866(.A(new_n894), .B1(new_n876), .B2(new_n881), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n891), .B1(new_n902), .B2(new_n903), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT39), .B1(new_n889), .B2(new_n867), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n738), .A2(new_n819), .A3(new_n880), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n819), .A2(new_n706), .A3(new_n674), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n873), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n880), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n890), .A2(new_n1074), .A3(new_n894), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n890), .A2(new_n1074), .A3(new_n894), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n893), .B2(new_n1067), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n899), .B1(new_n904), .B2(new_n732), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n880), .A2(new_n819), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n744), .B(new_n1076), .C1(new_n1078), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n748), .B1(new_n848), .B2(new_n249), .ZN(new_n1083));
  INV_X1    g0883(.A(G125), .ZN(new_n1084));
  INV_X1    g0884(.A(G132), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n271), .B1(new_n753), .B2(new_n1084), .C1(new_n778), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n769), .A2(G128), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n1048), .B2(new_n774), .C1(new_n220), .C2(new_n783), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT53), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n760), .B2(new_n251), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n761), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1086), .B(new_n1088), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n780), .A2(new_n828), .B1(new_n757), .B2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT109), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1055), .B1(G116), .B2(new_n765), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT110), .Z(new_n1097));
  OAI221_X1 g0897(.A(new_n350), .B1(new_n757), .B2(new_n583), .C1(new_n772), .C2(new_n753), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n780), .A2(new_n522), .B1(new_n768), .B2(new_n1017), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n1098), .A2(new_n834), .A3(new_n1099), .A4(new_n785), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1092), .A2(new_n1095), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1083), .B1(new_n750), .B2(new_n1101), .C1(new_n1102), .C2(new_n792), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1082), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n426), .A2(new_n1079), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n896), .A2(new_n639), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n876), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n880), .B1(new_n738), .B2(new_n819), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n1080), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n880), .B1(new_n819), .B2(new_n1079), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n1073), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1071), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT108), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1076), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1081), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1115), .B(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1113), .B(new_n1076), .C1(new_n1078), .C2(new_n1081), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1120), .A2(new_n693), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1104), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n902), .A2(new_n903), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n880), .B1(new_n813), .B2(new_n874), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1125), .A2(new_n1126), .B1(new_n636), .B2(new_n670), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n894), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1102), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n907), .A2(new_n908), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n899), .B1(new_n890), .B2(new_n909), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n670), .A2(new_n263), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n300), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n300), .A2(new_n1135), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n300), .A2(new_n1135), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1142), .B(KEYINPUT117), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1130), .A2(new_n1145), .A3(new_n1131), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1129), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1130), .A2(new_n1145), .A3(new_n1131), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n895), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1124), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1106), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1120), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n694), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1129), .A2(new_n1144), .A3(new_n1146), .A4(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1158), .B2(KEYINPUT57), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(G33), .A2(G41), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G50), .B(new_n1160), .C1(new_n831), .C2(new_n452), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT111), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n783), .A2(new_n385), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n760), .A2(new_n270), .B1(new_n753), .B2(new_n1017), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1163), .A2(new_n1164), .A3(G41), .A4(new_n799), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT112), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n778), .A2(new_n522), .B1(new_n337), .B2(new_n757), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n780), .A2(new_n583), .B1(new_n768), .B2(new_n429), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1166), .A2(new_n925), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1162), .B1(new_n1169), .B2(KEYINPUT58), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT113), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n780), .A2(new_n1085), .B1(new_n768), .B2(new_n1084), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n758), .A2(G137), .B1(G128), .B2(new_n765), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n760), .B2(new_n1093), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G150), .C2(new_n835), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT59), .Z(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT114), .ZN(new_n1177));
  OR2_X1    g0977(.A1(KEYINPUT115), .A2(G124), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(KEYINPUT115), .A2(G124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n754), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1160), .C1(new_n1048), .C2(new_n783), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1176), .B2(KEYINPUT114), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1177), .A2(new_n1182), .B1(KEYINPUT58), .B2(new_n1169), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n750), .B1(new_n1171), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT116), .Z(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n745), .C1(G50), .C2(new_n847), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1145), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n791), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n744), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1159), .A2(new_n1190), .ZN(G375));
  NAND2_X1  g0991(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n1152), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n978), .B(KEYINPUT119), .Z(new_n1195));
  NAND4_X1  g0995(.A1(new_n1115), .A2(new_n1194), .A3(new_n1116), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n881), .A2(new_n791), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n745), .B1(new_n847), .B2(G68), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n778), .A2(new_n1017), .B1(new_n757), .B2(new_n522), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n271), .B(new_n1199), .C1(G303), .C2(new_n754), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n835), .A2(new_n603), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n780), .A2(new_n429), .B1(new_n760), .B2(new_n583), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G294), .B2(new_n769), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n929), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n780), .A2(new_n1093), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1205), .B(new_n1163), .C1(G159), .C2(new_n761), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n769), .A2(G132), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n754), .A2(G128), .B1(G137), .B2(new_n765), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1208), .A3(new_n799), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n774), .A2(new_n220), .B1(new_n757), .B2(new_n251), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT121), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1198), .B1(new_n790), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT122), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1192), .A2(new_n744), .B1(new_n1197), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1196), .A2(new_n1216), .ZN(G381));
  OR3_X1    g1017(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G378), .A2(new_n1218), .A3(G381), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1065), .B(new_n950), .C1(new_n980), .C2(new_n998), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n1159), .A3(new_n1190), .A4(new_n1221), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n672), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1122), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G375), .C2(new_n1225), .ZN(G409));
  XNOR2_X1  g1026(.A(G393), .B(new_n807), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1034), .A2(new_n968), .A3(new_n967), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n978), .B1(new_n1228), .B2(new_n739), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n997), .B1(new_n1229), .B2(new_n744), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1065), .B1(new_n1230), .B2(new_n950), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1221), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(G390), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G393), .B(G396), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1220), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1159), .A2(G378), .A3(new_n1190), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1155), .A2(new_n1153), .A3(new_n1157), .A4(new_n1195), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1188), .B1(new_n1239), .B2(new_n744), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1122), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1244), .A3(new_n1122), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1237), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1113), .A2(new_n694), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1193), .A2(new_n1248), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1192), .A2(new_n1152), .A3(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1247), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1251), .B2(new_n1216), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(G384), .A3(new_n1216), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(KEYINPUT124), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1251), .A2(new_n1255), .A3(G384), .A4(new_n1216), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1246), .A2(new_n1223), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1223), .A4(new_n1257), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT62), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1223), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1224), .A2(G2897), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1252), .ZN(new_n1267));
  AND4_X1   g1067(.A1(new_n1256), .A2(new_n1266), .A3(new_n1267), .A4(new_n1264), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1236), .B1(new_n1262), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1232), .A2(new_n1274), .A3(new_n1235), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1232), .A2(new_n1235), .A3(new_n1277), .A4(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1263), .B2(new_n1269), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1260), .A2(new_n1281), .A3(new_n1261), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1258), .A2(new_n1281), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1273), .A2(new_n1284), .ZN(G405));
  NAND2_X1  g1085(.A1(G375), .A2(new_n1122), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(KEYINPUT127), .A3(new_n1237), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1287), .A2(new_n1236), .A3(new_n1257), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1236), .B1(new_n1287), .B2(new_n1257), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1286), .A2(new_n1237), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(KEYINPUT127), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1290), .B(new_n1292), .ZN(G402));
endmodule


