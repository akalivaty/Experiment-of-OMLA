//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n213), .A2(G50), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G200), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G222), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G223), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n248), .A2(G1698), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(new_n253), .B2(new_n248), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n258), .A2(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n264), .A2(G226), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n247), .B1(new_n260), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n260), .A2(new_n269), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(G190), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n216), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n217), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT67), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT8), .A2(G58), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT66), .B(G58), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(KEYINPUT8), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n275), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n274), .B1(new_n261), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n202), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n284), .A2(new_n290), .A3(KEYINPUT71), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT71), .B1(new_n284), .B2(new_n290), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n272), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n272), .B(new_n298), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n271), .A2(G169), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n284), .A2(new_n290), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n301), .A2(KEYINPUT68), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n271), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT68), .B1(new_n301), .B2(new_n302), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n201), .B1(new_n279), .B2(G68), .ZN(new_n310));
  INV_X1    g0110(.A(G159), .ZN(new_n311));
  INV_X1    g0111(.A(new_n282), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n310), .A2(new_n217), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n248), .B2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n241), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n309), .B1(new_n313), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT74), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n325), .A3(KEYINPUT7), .A4(new_n217), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n315), .ZN(new_n327));
  AOI21_X1  g0127(.A(G20), .B1(new_n317), .B2(new_n319), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n325), .B1(new_n328), .B2(KEYINPUT7), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT66), .A2(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT66), .A2(G58), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n201), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n217), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n312), .A2(new_n311), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n335), .A2(new_n309), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n275), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n309), .C1(new_n313), .C2(new_n322), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n324), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n289), .A2(new_n280), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n280), .B2(new_n286), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n268), .A2(new_n258), .A3(G274), .ZN(new_n344));
  INV_X1    g0144(.A(G232), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n263), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n248), .A2(G226), .A3(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G87), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n346), .B1(new_n350), .B2(new_n259), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G200), .B2(new_n351), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(new_n343), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n343), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n304), .B(new_n346), .C1(new_n259), .C2(new_n350), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI211_X1 g0165(.A(KEYINPUT18), .B(new_n365), .C1(new_n343), .C2(new_n341), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n341), .A2(new_n343), .ZN(new_n368));
  INV_X1    g0168(.A(new_n365), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n357), .A2(KEYINPUT75), .A3(new_n358), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n361), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(G226), .A2(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n345), .A2(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n248), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n259), .ZN(new_n379));
  INV_X1    g0179(.A(G238), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n344), .B1(new_n380), .B2(new_n263), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT13), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n258), .B1(new_n376), .B2(new_n377), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT13), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G190), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n277), .A2(G77), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n241), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n394));
  AOI22_X1  g0194(.A1(G68), .A2(new_n288), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT11), .B1(new_n391), .B2(new_n274), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n387), .A2(new_n247), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n398), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT72), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(KEYINPUT14), .C1(new_n387), .C2(new_n362), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n362), .B1(new_n384), .B2(new_n386), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT72), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n387), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n406), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n404), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n401), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n255), .A2(new_n380), .B1(new_n206), .B2(new_n248), .ZN(new_n412));
  OR3_X1    g0212(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n345), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT69), .B1(new_n250), .B2(new_n345), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n258), .ZN(new_n416));
  INV_X1    g0216(.A(G244), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n344), .B1(new_n263), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G190), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n286), .A2(new_n253), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n289), .B2(new_n253), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT8), .B(G58), .Z(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT15), .B(G87), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n276), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n274), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT70), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n427), .B(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n420), .B(new_n429), .C1(new_n247), .C2(new_n419), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n304), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n427), .B(KEYINPUT70), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n362), .B1(new_n416), .B2(new_n418), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n411), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n308), .A2(new_n373), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT25), .B1(new_n286), .B2(new_n206), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n261), .A2(G33), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n275), .A2(new_n285), .A3(new_n440), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n438), .A2(new_n439), .B1(new_n441), .B2(new_n206), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n317), .A2(new_n319), .A3(G257), .A4(G1698), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n317), .A2(new_n319), .A3(G250), .A4(new_n249), .ZN(new_n444));
  AND2_X1   g0244(.A1(KEYINPUT84), .A2(G294), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT84), .A2(G294), .ZN(new_n446));
  OAI21_X1  g0246(.A(G33), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n259), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n258), .A2(G274), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n267), .A2(G1), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(G264), .A3(new_n258), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n449), .A2(new_n352), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n449), .A2(new_n455), .A3(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n247), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n317), .A2(new_n319), .A3(new_n217), .A4(G87), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n248), .A2(new_n462), .A3(new_n217), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT23), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n217), .B2(G107), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n217), .A2(G33), .A3(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .A3(KEYINPUT24), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n464), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n461), .B2(new_n463), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n474), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n480), .A3(new_n474), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(new_n476), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  AOI221_X4 g0282(.A(new_n442), .B1(new_n457), .B2(new_n459), .C1(new_n482), .C2(new_n274), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n458), .A2(new_n362), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G179), .B2(new_n458), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n274), .ZN(new_n486));
  INV_X1    g0286(.A(new_n442), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n317), .A2(new_n319), .A3(G264), .A4(G1698), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT80), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n248), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n317), .A2(new_n319), .A3(G257), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n249), .B1(G303), .B2(new_n320), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n258), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n304), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n454), .A2(G270), .A3(new_n258), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n454), .A2(KEYINPUT79), .A3(G270), .A4(new_n258), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n455), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n286), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n273), .A2(new_n216), .B1(G20), .B2(new_n505), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n217), .C1(G33), .C2(new_n205), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(KEYINPUT20), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT20), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  OAI221_X1 g0311(.A(new_n506), .B1(new_n441), .B2(new_n505), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n498), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n497), .A2(new_n503), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n506), .B1(new_n441), .B2(new_n505), .ZN(new_n518));
  OAI21_X1  g0318(.A(G169), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n515), .B(KEYINPUT21), .C1(new_n516), .C2(new_n519), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(G190), .ZN(new_n525));
  INV_X1    g0325(.A(new_n512), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n247), .C2(new_n516), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n317), .A2(new_n319), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n317), .A2(new_n319), .A3(G244), .A4(new_n249), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n508), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n259), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n450), .A2(new_n454), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n454), .A2(new_n258), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(G257), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n362), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n205), .A3(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n217), .B1(new_n253), .B2(new_n312), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n206), .B1(new_n315), .B2(new_n321), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n274), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n285), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(new_n441), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n533), .A2(new_n536), .A3(new_n304), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G116), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n250), .B2(new_n380), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n255), .A2(new_n417), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n259), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n451), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n556), .A2(G250), .A3(new_n258), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n265), .A2(KEYINPUT76), .A3(new_n451), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT76), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n450), .B2(new_n556), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(new_n561), .A3(G190), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT78), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n555), .A2(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n555), .A2(new_n561), .A3(KEYINPUT78), .A4(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n248), .A2(new_n217), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n217), .B1(new_n377), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G87), .B2(new_n207), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n276), .B2(new_n205), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n274), .B1(new_n286), .B2(new_n425), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n547), .A2(G87), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n441), .A2(new_n425), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n574), .A2(KEYINPUT77), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT77), .B1(new_n574), .B2(new_n578), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n555), .A2(new_n561), .A3(G179), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n362), .B1(new_n555), .B2(new_n561), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n537), .A2(G200), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n533), .A2(new_n536), .A3(G190), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(new_n545), .A3(new_n548), .A4(new_n585), .ZN(new_n586));
  AND4_X1   g0386(.A1(new_n551), .A2(new_n577), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n489), .A2(new_n524), .A3(new_n527), .A4(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n437), .A2(new_n588), .ZN(G372));
  INV_X1    g0389(.A(new_n485), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT83), .B1(new_n472), .B2(KEYINPUT24), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n478), .A2(new_n477), .A3(new_n474), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n480), .A2(new_n464), .A3(new_n474), .A4(new_n471), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n480), .B1(new_n478), .B2(new_n474), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n275), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n590), .B1(new_n597), .B2(new_n442), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n524), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n566), .A2(new_n576), .A3(new_n562), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n586), .A2(new_n600), .A3(new_n551), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n483), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n574), .A2(new_n578), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n581), .B2(new_n582), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n600), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n551), .ZN(new_n608));
  INV_X1    g0408(.A(new_n551), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n577), .A3(new_n583), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n436), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n307), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n357), .A2(KEYINPUT75), .A3(new_n358), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT75), .B1(new_n357), .B2(new_n358), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n410), .A2(new_n402), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n401), .B2(new_n434), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n371), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n614), .B1(new_n621), .B2(new_n300), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n613), .A2(new_n622), .ZN(G369));
  INV_X1    g0423(.A(new_n524), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n261), .A2(new_n217), .A3(G13), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G213), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n526), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n524), .A2(new_n527), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G330), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n489), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n486), .B2(new_n487), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n639), .A2(new_n640), .B1(new_n598), .B2(new_n632), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n632), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n524), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n489), .B1(new_n488), .B2(new_n632), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(G399));
  NOR3_X1   g0446(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT86), .Z(new_n648));
  INV_X1    g0448(.A(new_n210), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n261), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n648), .A2(new_n651), .B1(new_n215), .B2(new_n650), .ZN(new_n652));
  XOR2_X1   g0452(.A(new_n652), .B(KEYINPUT28), .Z(new_n653));
  INV_X1    g0453(.A(new_n605), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n599), .B2(new_n602), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n643), .B1(new_n655), .B2(new_n611), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT29), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(KEYINPUT88), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n656), .B2(KEYINPUT29), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n607), .A2(new_n551), .ZN(new_n662));
  MUX2_X1   g0462(.A(new_n610), .B(new_n662), .S(KEYINPUT26), .Z(new_n663));
  AOI21_X1  g0463(.A(new_n643), .B1(new_n655), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT29), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n588), .A2(KEYINPUT31), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n449), .A2(new_n456), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n516), .B1(new_n455), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n304), .A3(new_n537), .A4(new_n565), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n498), .A2(new_n533), .A3(new_n536), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n669), .A2(new_n504), .A3(new_n555), .A4(new_n561), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n673), .A2(new_n674), .A3(new_n672), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n643), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT87), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n684), .B2(new_n676), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n632), .A2(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n667), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n666), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n653), .B1(new_n691), .B2(G1), .ZN(G364));
  AOI21_X1  g0492(.A(new_n216), .B1(G20), .B2(new_n362), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n217), .A2(new_n304), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G200), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n352), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT92), .B(G326), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n445), .A2(new_n446), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n352), .A2(G179), .A3(G200), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n217), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n700), .A2(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n697), .A2(G190), .A3(new_n247), .ZN(new_n708));
  INV_X1    g0508(.A(G322), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n320), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G190), .A2(G200), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n697), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(G311), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n698), .A2(G190), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT33), .B(G317), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n217), .A2(G179), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(G190), .A3(G200), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n715), .A2(new_n716), .B1(new_n719), .B2(G303), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n707), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n352), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(G283), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n717), .A2(new_n711), .ZN(new_n724));
  INV_X1    g0524(.A(G329), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n705), .A2(new_n706), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n721), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n704), .A2(new_n205), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n715), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n731), .B1(new_n206), .B2(new_n722), .C1(new_n241), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n724), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G159), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  INV_X1    g0536(.A(new_n279), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n248), .B1(new_n712), .B2(new_n253), .C1(new_n737), .C2(new_n708), .ZN(new_n738));
  INV_X1    g0538(.A(G87), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n700), .A2(new_n202), .B1(new_n718), .B2(new_n739), .ZN(new_n740));
  NOR4_X1   g0540(.A1(new_n733), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n696), .B1(new_n729), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n696), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n649), .A2(new_n320), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(G355), .B1(new_n505), .B2(new_n649), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n649), .A2(new_n248), .ZN(new_n750));
  INV_X1    g0550(.A(new_n215), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n751), .B2(G45), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n245), .A2(new_n267), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n747), .B1(new_n754), .B2(KEYINPUT89), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(KEYINPUT89), .B2(new_n754), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n217), .A2(G13), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n261), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n650), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n742), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT95), .ZN(new_n762));
  INV_X1    g0562(.A(new_n745), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n636), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n760), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n637), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n636), .A2(G330), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(G396));
  NOR2_X1   g0568(.A1(new_n434), .A2(new_n643), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n430), .B1(new_n429), .B2(new_n632), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n434), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n657), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n612), .A2(new_n771), .A3(new_n632), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(KEYINPUT98), .A3(new_n774), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n771), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(new_n690), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n690), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n778), .A2(new_n760), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(KEYINPUT99), .B2(new_n777), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n696), .A2(new_n743), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n765), .B1(new_n782), .B2(new_n253), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n723), .A2(new_n732), .B1(new_n700), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G107), .B2(new_n719), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n708), .A2(new_n788), .B1(new_n724), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n248), .B(new_n790), .C1(G116), .C2(new_n713), .ZN(new_n791));
  INV_X1    g0591(.A(new_n722), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n730), .B1(G87), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n248), .B1(new_n724), .B2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n704), .A2(new_n737), .B1(new_n718), .B2(new_n202), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G68), .C2(new_n792), .ZN(new_n798));
  INV_X1    g0598(.A(new_n708), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT97), .B(G143), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(new_n801), .B1(new_n713), .B2(G159), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n699), .A2(G137), .ZN(new_n803));
  INV_X1    g0603(.A(G150), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n732), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n806), .B2(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT34), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n794), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n784), .B1(new_n810), .B2(new_n696), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n771), .B2(new_n744), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n781), .A2(new_n812), .ZN(G384));
  INV_X1    g0613(.A(new_n542), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT35), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(KEYINPUT35), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n815), .A2(G116), .A3(new_n218), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT36), .Z(new_n818));
  NAND3_X1  g0618(.A1(new_n215), .A2(G77), .A3(new_n333), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n240), .B(KEYINPUT100), .Z(new_n820));
  AOI211_X1 g0620(.A(new_n261), .B(G13), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT102), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n769), .B1(new_n656), .B2(new_n771), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n401), .A2(new_n410), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n402), .A2(new_n643), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n401), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n618), .A2(new_n828), .A3(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n411), .A2(KEYINPUT101), .A3(new_n826), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n823), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n769), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n774), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n833), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT102), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n368), .A2(new_n369), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n368), .A2(new_n631), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n355), .ZN(new_n844));
  INV_X1    g0644(.A(new_n338), .ZN(new_n845));
  INV_X1    g0645(.A(new_n313), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT16), .B1(new_n330), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n343), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n369), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n631), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n355), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  INV_X1    g0652(.A(new_n850), .ZN(new_n853));
  AOI221_X4 g0653(.A(new_n840), .B1(new_n844), .B2(new_n852), .C1(new_n373), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n373), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n844), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT103), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n850), .B1(new_n617), .B2(new_n371), .ZN(new_n859));
  INV_X1    g0659(.A(new_n856), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n840), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n855), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n839), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  INV_X1    g0666(.A(new_n842), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n357), .A2(new_n868), .A3(new_n358), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n371), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n868), .B1(new_n357), .B2(new_n358), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n841), .A2(new_n842), .A3(new_n355), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n844), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n866), .B1(new_n854), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n863), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n618), .A2(new_n643), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n371), .A2(new_n631), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT105), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n858), .A2(new_n864), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n834), .A3(new_n838), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n880), .A4(new_n881), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n659), .A2(new_n436), .A3(new_n661), .A4(new_n665), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n622), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n888), .B(new_n890), .Z(new_n891));
  NAND2_X1  g0691(.A1(new_n677), .A2(new_n680), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n668), .A2(new_n682), .B1(new_n892), .B2(new_n687), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n837), .A3(new_n771), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n858), .B2(new_n864), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT40), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n893), .A2(new_n833), .A3(new_n898), .A4(new_n772), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n872), .A2(new_n875), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n840), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n863), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n437), .B2(new_n893), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n897), .A2(new_n436), .A3(new_n894), .A4(new_n903), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(G330), .A3(new_n906), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n891), .A2(new_n907), .B1(new_n261), .B2(new_n757), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT106), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n891), .A2(new_n907), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(KEYINPUT106), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n822), .B1(new_n911), .B2(new_n912), .ZN(G367));
  OAI21_X1  g0713(.A(new_n746), .B1(new_n210), .B2(new_n425), .ZN(new_n914));
  INV_X1    g0714(.A(new_n750), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n235), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n760), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n704), .A2(new_n241), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G150), .B2(new_n799), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT113), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n732), .A2(new_n311), .B1(new_n737), .B2(new_n718), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n700), .A2(new_n800), .B1(new_n253), .B2(new_n722), .ZN(new_n922));
  XOR2_X1   g0722(.A(KEYINPUT114), .B(G137), .Z(new_n923));
  OAI221_X1 g0723(.A(new_n248), .B1(new_n712), .B2(new_n202), .C1(new_n724), .C2(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n799), .A2(G303), .B1(new_n713), .B2(G283), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n206), .B2(new_n704), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n702), .A2(new_n732), .B1(new_n700), .B2(new_n789), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n718), .A2(new_n505), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT46), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(G317), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n320), .B1(new_n724), .B2(new_n932), .C1(new_n205), .C2(new_n722), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT112), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n920), .A2(new_n925), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT47), .ZN(new_n936));
  INV_X1    g0736(.A(new_n696), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(KEYINPUT47), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n917), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n632), .A2(new_n576), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n654), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n607), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n942), .B2(new_n763), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n643), .A2(new_n549), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n551), .A3(new_n586), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n609), .A2(new_n643), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n645), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n944), .B1(new_n645), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n645), .A2(new_n949), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n645), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n638), .A3(new_n641), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT110), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n952), .A2(new_n957), .A3(new_n642), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n644), .A2(new_n489), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n641), .B2(new_n644), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(KEYINPUT111), .B2(new_n637), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n637), .B(KEYINPUT111), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n691), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n691), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n650), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n759), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT107), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(KEYINPUT108), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n965), .A2(new_n948), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT42), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n551), .B1(new_n598), .B2(new_n946), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n632), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n978), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n977), .A2(KEYINPUT108), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT109), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n642), .A2(new_n948), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(KEYINPUT109), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n987), .B(new_n988), .C1(new_n985), .C2(new_n986), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n943), .B1(new_n974), .B2(new_n993), .ZN(G387));
  NAND2_X1  g0794(.A1(new_n969), .A2(new_n759), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n750), .B1(new_n232), .B2(new_n267), .ZN(new_n996));
  INV_X1    g0796(.A(new_n748), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n648), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n267), .B1(new_n241), .B2(new_n253), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n423), .A2(new_n202), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n648), .B(new_n1001), .C1(KEYINPUT50), .C2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n998), .A2(new_n1002), .B1(new_n206), .B2(new_n649), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n760), .B1(new_n1003), .B2(new_n747), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n799), .A2(G317), .B1(new_n713), .B2(G303), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n700), .B2(new_n709), .C1(new_n789), .C2(new_n732), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n723), .B2(new_n704), .C1(new_n702), .C2(new_n718), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n320), .B1(new_n724), .B2(new_n701), .C1(new_n505), .C2(new_n722), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT49), .B2(new_n1011), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n712), .A2(new_n241), .B1(new_n724), .B2(new_n804), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n320), .B(new_n1016), .C1(G50), .C2(new_n799), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n704), .A2(new_n425), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n792), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n699), .A2(G159), .B1(new_n719), .B2(G77), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n715), .A2(new_n280), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1004), .B1(new_n1023), .B2(new_n696), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n641), .B2(new_n763), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n970), .A2(new_n650), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n691), .A2(new_n969), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n995), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(G393));
  NAND3_X1  g0828(.A1(new_n959), .A2(new_n759), .A3(new_n963), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n704), .A2(new_n253), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n713), .A2(new_n423), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n732), .B2(new_n202), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1032), .B2(KEYINPUT115), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(KEYINPUT115), .B2(new_n1032), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT116), .Z(new_n1035));
  OAI22_X1  g0835(.A1(new_n700), .A2(new_n804), .B1(new_n311), .B2(new_n708), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n248), .B1(new_n724), .B2(new_n800), .C1(new_n739), .C2(new_n722), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G68), .B2(new_n719), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G317), .A2(new_n699), .B1(new_n799), .B2(G311), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n320), .B1(new_n724), .B2(new_n709), .C1(new_n788), .C2(new_n712), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n732), .A2(new_n785), .B1(new_n722), .B2(new_n206), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n704), .A2(new_n505), .B1(new_n718), .B2(new_n723), .ZN(new_n1045));
  OR4_X1    g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n937), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n239), .A2(new_n915), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n747), .B1(G97), .B2(new_n649), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n765), .B(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n763), .B2(new_n949), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1029), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT117), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n959), .A2(new_n963), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n970), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n650), .B(new_n1056), .C1(new_n964), .C2(new_n970), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n1057), .ZN(G390));
  NAND2_X1  g0858(.A1(new_n836), .A2(new_n837), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n879), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n878), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT39), .B1(new_n901), .B2(new_n863), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n879), .B(KEYINPUT118), .Z(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n854), .B2(new_n876), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n770), .A2(new_n434), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n769), .B1(new_n664), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(new_n833), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n689), .A2(new_n771), .A3(new_n837), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1064), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n893), .A2(new_n833), .A3(new_n667), .A4(new_n772), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n877), .A2(new_n878), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n1070), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1076), .A3(new_n759), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n782), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n760), .B1(new_n1078), .B2(new_n280), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n712), .A2(new_n205), .B1(new_n724), .B2(new_n788), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G116), .B2(new_n799), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1030), .B1(G68), .B2(new_n792), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n715), .A2(G107), .B1(new_n699), .B2(G283), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n320), .B1(new_n718), .B2(new_n739), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT120), .Z(new_n1086));
  NAND2_X1  g0886(.A1(new_n719), .A2(G150), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT53), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n704), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n923), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G159), .A2(new_n1089), .B1(new_n715), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n708), .A2(new_n795), .B1(new_n724), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n248), .B1(new_n712), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n699), .A2(G128), .B1(new_n792), .B2(G50), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1091), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1084), .A2(new_n1086), .B1(new_n1088), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1099), .B2(new_n696), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n744), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1077), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n894), .A2(new_n436), .A3(G330), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n889), .A2(new_n622), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n837), .B1(new_n689), .B2(new_n771), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n836), .B1(new_n1108), .B2(new_n1074), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n893), .A2(new_n667), .A3(new_n772), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1072), .B(new_n1068), .C1(new_n1110), .C2(new_n837), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(KEYINPUT119), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1073), .A2(new_n1112), .A3(new_n1076), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n650), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1104), .A2(new_n1105), .B1(new_n1116), .B2(new_n1118), .ZN(G378));
  AOI21_X1  g0919(.A(new_n667), .B1(new_n899), .B2(new_n902), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n896), .B2(KEYINPUT40), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n293), .A2(new_n631), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n308), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n1120), .C1(new_n896), .C2(KEYINPUT40), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n888), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n883), .A3(new_n887), .A4(new_n1128), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n759), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n760), .B1(new_n1078), .B2(G50), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n248), .A2(G41), .ZN(new_n1134));
  AOI211_X1 g0934(.A(G50), .B(new_n1134), .C1(new_n316), .C2(new_n266), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1134), .B1(new_n723), .B2(new_n724), .C1(new_n425), .C2(new_n712), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n918), .B(new_n1136), .C1(G77), .C2(new_n719), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n699), .A2(G116), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n715), .A2(G97), .B1(new_n792), .B2(new_n279), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n708), .A2(new_n206), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT122), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT58), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(KEYINPUT123), .A2(G124), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(KEYINPUT123), .A2(G124), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n734), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1147), .A2(new_n316), .A3(new_n266), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1092), .A2(new_n700), .B1(new_n732), .B2(new_n795), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n799), .A2(G128), .B1(new_n713), .B2(G137), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n718), .B2(new_n1094), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G150), .C2(new_n1089), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT59), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1148), .B1(new_n311), .B2(new_n722), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1152), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1144), .B1(new_n1143), .B2(new_n1142), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1133), .B1(new_n1157), .B2(new_n696), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1125), .B2(new_n744), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1132), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1107), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1117), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1130), .A2(new_n1162), .A3(new_n1131), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1130), .A2(KEYINPUT57), .A3(new_n1162), .A4(new_n1131), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n650), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1165), .B2(new_n1167), .ZN(G375));
  AND2_X1   g0968(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(new_n758), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n833), .A2(new_n743), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n765), .B1(new_n782), .B2(new_n241), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n248), .B1(new_n734), .B2(G303), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n206), .B2(new_n712), .C1(new_n723), .C2(new_n708), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1018), .B(new_n1174), .C1(G77), .C2(new_n792), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n505), .A2(new_n732), .B1(new_n700), .B2(new_n788), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G97), .B2(new_n719), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n719), .A2(G159), .B1(new_n734), .B2(G128), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT124), .Z(new_n1179));
  OAI22_X1  g0979(.A1(new_n795), .A2(new_n700), .B1(new_n732), .B2(new_n1094), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n248), .B1(new_n712), .B2(new_n804), .C1(new_n708), .C2(new_n923), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n704), .A2(new_n202), .B1(new_n737), .B2(new_n722), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1175), .A2(new_n1177), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1171), .B(new_n1172), .C1(new_n937), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1170), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n972), .B1(new_n1169), .B2(new_n1107), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G381));
  NOR4_X1   g0990(.A1(G390), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n974), .A2(new_n993), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1191), .A2(new_n943), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1132), .A2(new_n1159), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1166), .A2(new_n650), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1077), .B(new_n1102), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1193), .A2(new_n1197), .A3(new_n1189), .A4(new_n1199), .ZN(G407));
  INV_X1    g1000(.A(G343), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(G213), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT125), .Z(new_n1203));
  NAND3_X1  g1003(.A1(new_n1197), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(G407), .A2(G213), .A3(new_n1204), .ZN(G409));
  OAI211_X1 g1005(.A(G378), .B(new_n1160), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1163), .A2(new_n972), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1199), .B1(new_n1194), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1202), .ZN(new_n1210));
  INV_X1    g1010(.A(G384), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1212), .A2(new_n650), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1169), .A2(new_n1107), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n1112), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1211), .B1(new_n1217), .B2(new_n1186), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1186), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(G384), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1218), .A2(new_n1220), .B1(G2897), .B2(new_n1203), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1201), .A2(G213), .A3(G2897), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1218), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1210), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1209), .A2(new_n1202), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT63), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1203), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(KEYINPUT63), .A3(new_n1226), .ZN(new_n1231));
  XOR2_X1   g1031(.A(G393), .B(G396), .Z(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G390), .ZN(new_n1234));
  AND2_X1   g1034(.A1(G387), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G387), .A2(new_n1234), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1192), .A2(new_n943), .A3(G390), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1234), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1232), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(KEYINPUT61), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1224), .A2(new_n1229), .A3(new_n1231), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1223), .A2(new_n1221), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1227), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1230), .A2(KEYINPUT62), .A3(new_n1226), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1243), .B1(new_n1250), .B2(new_n1251), .ZN(G405));
  OAI211_X1 g1052(.A(new_n1206), .B(new_n1225), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G375), .A2(new_n1199), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1225), .B1(new_n1255), .B2(new_n1206), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1251), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(KEYINPUT127), .B(new_n1251), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1206), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1196), .A2(new_n650), .A3(new_n1166), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1198), .B1(new_n1262), .B2(new_n1160), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1226), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1241), .A3(new_n1253), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1241), .A3(new_n1267), .A4(new_n1253), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1259), .A2(new_n1260), .B1(new_n1266), .B2(new_n1268), .ZN(G402));
endmodule


