//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT1), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(KEYINPUT70), .A3(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n208), .ZN(new_n215));
  OR2_X1    g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(G134gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT69), .B(G127gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT24), .A3(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n222), .A2(KEYINPUT24), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT23), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n223), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n226), .B2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n234), .B(new_n235), .C1(G169gat), .C2(G176gat), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n237), .A3(KEYINPUT66), .ZN(new_n238));
  AND2_X1   g037(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT23), .B(new_n230), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n223), .A3(new_n224), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n225), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n224), .A3(new_n227), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(new_n243), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n238), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n231), .A2(KEYINPUT26), .A3(new_n226), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n222), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n254));
  AOI21_X1  g053(.A(G190gat), .B1(new_n254), .B2(KEYINPUT27), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(new_n261), .A3(new_n257), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT27), .B(G183gat), .Z(new_n264));
  OR3_X1    g063(.A1(new_n264), .A2(new_n260), .A3(G190gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n253), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n220), .B1(new_n248), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n252), .ZN(new_n269));
  MUX2_X1   g068(.A(G127gat), .B(new_n218), .S(G134gat), .Z(new_n270));
  AOI22_X1  g069(.A1(new_n212), .A2(new_n213), .B1(new_n270), .B2(new_n215), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n238), .A2(new_n244), .A3(new_n247), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G227gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n203), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n267), .A2(KEYINPUT34), .A3(new_n279), .A4(new_n273), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  AOI21_X1  g084(.A(new_n279), .B1(new_n267), .B2(new_n273), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(KEYINPUT33), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT32), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n271), .B1(new_n269), .B2(new_n272), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n277), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  INV_X1    g093(.A(new_n285), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n293), .B(KEYINPUT32), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n282), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n294), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n285), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n281), .A3(new_n296), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n302), .A2(KEYINPUT71), .A3(new_n281), .A4(new_n296), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G85gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315));
  OR2_X1    g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(KEYINPUT2), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n317), .B(new_n316), .C1(new_n321), .C2(KEYINPUT2), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n214), .A2(new_n323), .A3(new_n324), .A4(new_n219), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n271), .A2(KEYINPUT76), .A3(new_n324), .A4(new_n323), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n214), .A2(new_n323), .A3(new_n219), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(new_n322), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n220), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n220), .A2(new_n334), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n333), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n220), .A2(KEYINPUT77), .A3(new_n334), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(KEYINPUT5), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n329), .A2(new_n330), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n333), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n314), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n314), .A3(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT6), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n352), .B2(KEYINPUT6), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(G197gat), .ZN(new_n367));
  INV_X1    g166(.A(G204gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n365), .B(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n362), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n334), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(G228gat), .B2(G233gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(KEYINPUT29), .B2(new_n335), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n378), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G50gat), .ZN(new_n383));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(KEYINPUT80), .B2(G22gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(G22gat), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT35), .ZN(new_n389));
  INV_X1    g188(.A(new_n387), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n379), .A2(new_n380), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n269), .A2(new_n272), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT73), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G226gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n276), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n269), .A2(KEYINPUT73), .A3(new_n272), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n372), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(KEYINPUT29), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n393), .A2(new_n396), .A3(new_n276), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n395), .A2(new_n398), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(new_n400), .ZN(new_n407));
  XOR2_X1   g206(.A(G8gat), .B(G36gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G64gat), .ZN(new_n409));
  INV_X1    g208(.A(G92gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n407), .A2(new_n416), .A3(KEYINPUT30), .A4(new_n412), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n412), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n403), .B(new_n411), .C1(new_n406), .C2(new_n400), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n361), .A2(new_n392), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n202), .B1(new_n309), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n352), .A2(KEYINPUT6), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n356), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n415), .A3(new_n417), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n388), .A2(new_n391), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n298), .A2(new_n303), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT35), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n304), .A2(new_n306), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT84), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n304), .A2(new_n306), .A3(new_n305), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(KEYINPUT83), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n346), .A2(new_n314), .A3(new_n351), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n352), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n439), .A2(new_n358), .B1(new_n441), .B2(new_n355), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n442), .A2(new_n428), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n444), .A3(KEYINPUT85), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n434), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n405), .A2(new_n401), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n400), .C1(new_n448), .C2(new_n404), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n399), .A2(new_n372), .A3(new_n402), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT82), .B1(new_n406), .B2(new_n372), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT37), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n412), .B1(new_n407), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n407), .A2(new_n454), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n457), .A2(KEYINPUT38), .A3(new_n455), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n413), .B(new_n442), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n431), .ZN(new_n460));
  INV_X1    g259(.A(new_n342), .ZN(new_n461));
  INV_X1    g260(.A(new_n344), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n333), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n347), .A2(new_n343), .A3(new_n348), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT39), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n314), .B1(new_n464), .B2(KEYINPUT39), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(new_n428), .A3(new_n353), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n459), .A2(new_n460), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n430), .A2(new_n431), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n304), .A2(new_n306), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n298), .A2(KEYINPUT36), .A3(new_n303), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n446), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G190gat), .B(G218gat), .Z(new_n482));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT15), .B(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n487), .A2(new_n488), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(G50gat), .ZN(new_n496));
  INV_X1    g295(.A(G50gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(G43gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n492), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(KEYINPUT87), .A2(KEYINPUT17), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n501), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(G85gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(KEYINPUT8), .A2(new_n510), .B1(new_n511), .B2(new_n410), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n511), .B2(new_n410), .ZN(new_n514));
  NAND3_X1  g313(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G99gat), .B(G106gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n509), .A2(new_n518), .B1(KEYINPUT41), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n517), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n516), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n501), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n482), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n482), .A3(new_n523), .ZN(new_n526));
  XOR2_X1   g325(.A(G134gat), .B(G162gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT94), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n519), .A2(KEYINPUT41), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  AND4_X1   g329(.A1(KEYINPUT95), .A2(new_n525), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n520), .A2(new_n532), .A3(new_n482), .A4(new_n523), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n525), .A2(new_n526), .B1(new_n533), .B2(new_n530), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G15gat), .A2(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(G15gat), .A2(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G15gat), .ZN(new_n550));
  INV_X1    g349(.A(G22gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT88), .B1(new_n552), .B2(new_n545), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT16), .ZN(new_n554));
  OAI22_X1  g353(.A1(new_n549), .A2(new_n553), .B1(new_n554), .B2(G1gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(G1gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n545), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n556), .A2(new_n558), .B1(KEYINPUT16), .B2(new_n557), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n562));
  OAI21_X1  g361(.A(G8gat), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G8gat), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n555), .B(new_n559), .C1(KEYINPUT89), .C2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G183gat), .ZN(new_n571));
  AND2_X1   g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574));
  INV_X1    g373(.A(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n573), .A2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n544), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n543), .A3(new_n578), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n535), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT11), .B(G169gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(G113gat), .B(G141gat), .Z(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT86), .Z(new_n590));
  OAI21_X1  g389(.A(new_n501), .B1(new_n564), .B2(new_n567), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n555), .A2(new_n559), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(G8gat), .C1(new_n562), .C2(new_n561), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n566), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT90), .A3(new_n501), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n568), .B1(new_n507), .B2(new_n508), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n568), .A2(new_n502), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT90), .B1(new_n596), .B2(new_n501), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n592), .B(new_n502), .C1(new_n595), .C2(new_n566), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n599), .B(KEYINPUT13), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n601), .B2(new_n607), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n590), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n601), .A2(new_n607), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n618), .A3(new_n613), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n589), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n230), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G204gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627));
  INV_X1    g426(.A(new_n539), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n538), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n517), .A2(KEYINPUT96), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n518), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n540), .A2(new_n522), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G230gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n276), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n627), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n627), .A3(new_n636), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n540), .A2(new_n522), .A3(KEYINPUT10), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n636), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n626), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  INV_X1    g446(.A(new_n626), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n647), .A2(new_n648), .A3(new_n644), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n623), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n640), .A2(new_n626), .A3(new_n645), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n648), .B1(new_n647), .B2(new_n644), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT98), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n622), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n481), .A2(new_n584), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n427), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n557), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n429), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n554), .A2(new_n565), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT42), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(KEYINPUT42), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n664), .B(new_n665), .C1(new_n565), .C2(new_n660), .ZN(G1325gat));
  OAI21_X1  g465(.A(new_n550), .B1(new_n657), .B2(new_n309), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT99), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n657), .A2(new_n550), .A3(new_n479), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n657), .A2(new_n460), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n481), .A2(new_n535), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n581), .A2(new_n583), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n656), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n485), .A3(new_n426), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  NAND2_X1  g480(.A1(KEYINPUT101), .A2(KEYINPUT44), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT101), .A2(KEYINPUT44), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n481), .B2(new_n535), .ZN(new_n687));
  INV_X1    g486(.A(new_n535), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n688), .B(new_n682), .C1(new_n446), .C2(new_n480), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n677), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n427), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n681), .A2(new_n693), .ZN(G1328gat));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n486), .A3(new_n428), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n692), .B2(new_n429), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n692), .B2(new_n479), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n688), .B1(new_n446), .B2(new_n480), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n700), .A2(new_n495), .A3(new_n438), .A4(new_n691), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT103), .Z(new_n702));
  AOI21_X1  g501(.A(KEYINPUT102), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1330gat));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n431), .A3(new_n691), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G50gat), .ZN(new_n707));
  NOR4_X1   g506(.A1(new_n674), .A2(G50gat), .A3(new_n460), .A4(new_n677), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n711), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AND4_X1   g517(.A1(new_n713), .A2(new_n707), .A3(new_n717), .A4(new_n714), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n712), .B1(new_n718), .B2(new_n719), .ZN(G1331gat));
  NAND3_X1  g519(.A1(new_n584), .A2(new_n622), .A3(new_n655), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT106), .Z(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n481), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n426), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n481), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n428), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  INV_X1    g532(.A(G71gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n723), .A2(new_n734), .A3(new_n438), .ZN(new_n735));
  OAI21_X1  g534(.A(G71gat), .B1(new_n726), .B2(new_n479), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n735), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n431), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  INV_X1    g544(.A(new_n687), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n700), .A2(new_n683), .ZN(new_n747));
  INV_X1    g546(.A(new_n622), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n675), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n746), .A2(new_n655), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n427), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n481), .A2(new_n535), .A3(new_n749), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n654), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n511), .A3(new_n426), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n757), .ZN(G1336gat));
  NOR2_X1   g557(.A1(new_n728), .A2(G92gat), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT109), .B1(new_n754), .B2(new_n755), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT51), .B1(new_n700), .B2(new_n749), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n655), .B(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G92gat), .B1(new_n750), .B2(new_n429), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT110), .B1(new_n766), .B2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n768), .B(new_n769), .C1(new_n764), .C2(new_n765), .ZN(new_n770));
  AND4_X1   g569(.A1(KEYINPUT51), .A2(new_n481), .A3(new_n535), .A4(new_n749), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n655), .B(new_n759), .C1(new_n771), .C2(new_n761), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n755), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n655), .A4(new_n759), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(new_n728), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n690), .A2(new_n655), .A3(new_n780), .A4(new_n749), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(G92gat), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n777), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n777), .B2(new_n782), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n767), .A2(new_n770), .B1(new_n783), .B2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n750), .A2(new_n786), .A3(new_n479), .ZN(new_n787));
  AOI21_X1  g586(.A(G99gat), .B1(new_n756), .B2(new_n438), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1338gat));
  OR2_X1    g588(.A1(new_n750), .A2(new_n460), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n460), .A2(new_n654), .A3(G106gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(G106gat), .B1(new_n775), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n760), .A2(new_n763), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(new_n791), .B1(new_n790), .B2(G106gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n642), .A2(new_n643), .ZN(new_n799));
  INV_X1    g598(.A(new_n636), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n644), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT54), .B(new_n636), .C1(new_n642), .C2(new_n643), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n626), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n799), .A2(new_n806), .A3(new_n800), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(KEYINPUT115), .A3(new_n648), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n802), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n649), .B1(new_n809), .B2(KEYINPUT55), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n810), .B(KEYINPUT116), .C1(KEYINPUT55), .C2(new_n809), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n801), .A2(new_n644), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n804), .A2(new_n803), .A3(new_n626), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n807), .B2(new_n648), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n651), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n809), .A2(KEYINPUT55), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n811), .B(new_n820), .C1(new_n621), .C2(new_n615), .ZN(new_n821));
  INV_X1    g620(.A(new_n588), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n605), .A2(new_n606), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n599), .B1(new_n598), .B2(new_n600), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n620), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n655), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n535), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n535), .A2(new_n811), .A3(new_n820), .A4(new_n826), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n676), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n584), .A2(new_n622), .A3(new_n654), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n427), .A3(new_n780), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n309), .A2(new_n431), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n622), .ZN(new_n837));
  INV_X1    g636(.A(new_n433), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n748), .A2(new_n206), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n836), .B2(new_n654), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n655), .A2(new_n204), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n839), .B2(new_n843), .ZN(G1341gat));
  NOR3_X1   g643(.A1(new_n836), .A2(new_n218), .A3(new_n676), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n834), .A2(new_n675), .A3(new_n838), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n218), .B2(new_n846), .ZN(G1342gat));
  NOR3_X1   g646(.A1(new_n833), .A2(new_n427), .A3(new_n433), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n429), .A2(new_n535), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT117), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n217), .A3(new_n850), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT56), .Z(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n836), .B2(new_n688), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1343gat));
  AOI21_X1  g653(.A(new_n460), .B1(new_n830), .B2(new_n831), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n479), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n427), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n728), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT118), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n584), .A2(new_n622), .A3(new_n654), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n809), .B2(KEYINPUT55), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n816), .A2(KEYINPUT119), .A3(new_n817), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n810), .B(new_n866), .C1(new_n615), .C2(new_n621), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n535), .B1(new_n867), .B2(new_n827), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n676), .B1(new_n868), .B2(new_n829), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT120), .B(new_n676), .C1(new_n868), .C2(new_n829), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n460), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n857), .B(new_n861), .C1(new_n873), .C2(new_n856), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n622), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n855), .A2(new_n859), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n728), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n622), .A2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(new_n876), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n877), .A2(new_n728), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(KEYINPUT122), .A3(new_n879), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n878), .B2(new_n880), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  INV_X1    g686(.A(new_n861), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n870), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n831), .A3(new_n872), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n431), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n891), .B2(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n892), .B2(new_n857), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n748), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n886), .B1(new_n895), .B2(G141gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n881), .B1(new_n896), .B2(new_n876), .ZN(G1344gat));
  INV_X1    g696(.A(G148gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n898), .A3(new_n655), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n892), .A2(new_n887), .A3(new_n857), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n654), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n898), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n818), .A2(new_n819), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n535), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n535), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n908), .A2(new_n826), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n676), .B1(new_n911), .B2(new_n868), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT57), .B(new_n460), .C1(new_n912), .C2(new_n831), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n855), .A2(new_n856), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n905), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n855), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n915), .A2(new_n655), .A3(new_n861), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n904), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n899), .B1(new_n903), .B2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(G155gat), .B1(new_n882), .B2(new_n675), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n901), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n675), .A2(G155gat), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT125), .Z(new_n923));
  AOI21_X1  g722(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(G1346gat));
  INV_X1    g723(.A(G162gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n877), .A2(new_n925), .A3(new_n850), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n688), .B1(new_n900), .B2(new_n901), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n728), .A2(new_n426), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n832), .A2(new_n838), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n930), .B(new_n748), .C1(new_n240), .C2(new_n239), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n429), .A2(new_n426), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n832), .A2(new_n835), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n622), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1348gat));
  AOI21_X1  g734(.A(G176gat), .B1(new_n930), .B2(new_n655), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n933), .A2(new_n230), .A3(new_n654), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  NOR2_X1   g737(.A1(new_n676), .A2(new_n264), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G183gat), .B1(new_n933), .B2(new_n676), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT126), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n945));
  OAI221_X1 g744(.A(G190gat), .B1(KEYINPUT127), .B2(new_n945), .C1(new_n933), .C2(new_n688), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n535), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(G190gat), .B2(new_n949), .ZN(G1351gat));
  AND2_X1   g749(.A1(new_n855), .A2(new_n929), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n479), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n367), .A3(new_n748), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n915), .A2(new_n916), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n932), .A2(new_n479), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n748), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n957), .B2(new_n367), .ZN(G1352gat));
  NOR3_X1   g757(.A1(new_n952), .A2(G204gat), .A3(new_n654), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n955), .A2(new_n655), .A3(new_n956), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n368), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n953), .A2(new_n575), .A3(new_n675), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n915), .A2(new_n675), .A3(new_n916), .A4(new_n956), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n535), .A3(new_n956), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G218gat), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n952), .A2(G218gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n688), .B2(new_n970), .ZN(G1355gat));
endmodule


