//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .A3(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(G146), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n198), .B2(G119), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n200), .A2(G128), .B1(KEYINPUT78), .B2(KEYINPUT23), .ZN(new_n213));
  INV_X1    g027(.A(new_n211), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT79), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n216), .B2(new_n199), .ZN(new_n217));
  INV_X1    g031(.A(G110), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n205), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n197), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n210), .A2(new_n208), .A3(new_n211), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT79), .B1(new_n213), .B2(new_n214), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n199), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n218), .A3(new_n206), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n204), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT81), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT16), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n193), .A3(G125), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n196), .B2(new_n228), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n192), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n202), .A2(new_n203), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n218), .B1(new_n224), .B2(new_n206), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT80), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n212), .A2(new_n215), .B1(G119), .B2(new_n198), .ZN(new_n239));
  OAI21_X1  g053(.A(G110), .B1(new_n239), .B2(new_n207), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n232), .B2(new_n192), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n221), .A2(new_n227), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G137), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n245), .B(new_n247), .Z(new_n248));
  OAI21_X1  g062(.A(new_n187), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n225), .A2(new_n220), .A3(new_n204), .ZN(new_n250));
  INV_X1    g064(.A(new_n197), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n220), .B1(new_n225), .B2(new_n204), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n242), .B1(new_n240), .B2(new_n241), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n248), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(KEYINPUT82), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n249), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n244), .A2(new_n248), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT76), .B(G902), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G234), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G902), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n244), .B2(new_n248), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n227), .A2(new_n250), .A3(new_n251), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n238), .A2(new_n243), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n187), .B(new_n248), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT82), .B1(new_n256), .B2(new_n257), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n267), .B(KEYINPUT25), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n263), .B(KEYINPUT77), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n265), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT71), .B(G237), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(G210), .A3(new_n246), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT73), .Z(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G101), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n283), .B(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G113), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT2), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G113), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT66), .A2(G116), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(G119), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n200), .A2(G116), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n289), .A2(new_n291), .B1(G116), .B2(new_n200), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT67), .B1(new_n301), .B2(new_n297), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n298), .A3(new_n292), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT68), .A3(new_n300), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n231), .B2(G143), .ZN(new_n314));
  INV_X1    g128(.A(G143), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT65), .A3(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(G146), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT0), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n198), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT64), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n315), .B2(G146), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n317), .A2(new_n319), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n198), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n231), .A2(G143), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n325), .B(new_n326), .C1(new_n327), .C2(new_n318), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT11), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(G137), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G131), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n332), .A2(new_n334), .A3(new_n338), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT1), .ZN(new_n342));
  OAI21_X1  g156(.A(G128), .B1(new_n318), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n327), .B2(new_n318), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n317), .A2(new_n319), .A3(new_n323), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n331), .A2(G137), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n333), .A2(G134), .ZN(new_n349));
  OAI21_X1  g163(.A(G131), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n350), .A3(KEYINPUT69), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n347), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n306), .A2(new_n312), .A3(new_n341), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT70), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n306), .A2(new_n312), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n344), .A2(new_n346), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n341), .B1(new_n360), .B2(new_n351), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n344), .A2(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(new_n354), .B1(new_n329), .B2(new_n340), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(KEYINPUT70), .A3(new_n306), .A4(new_n312), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT28), .ZN(new_n367));
  INV_X1    g181(.A(new_n356), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT28), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n287), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n358), .A2(new_n373), .A3(new_n365), .A4(new_n287), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n341), .A2(new_n355), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(KEYINPUT30), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n361), .A2(KEYINPUT30), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n359), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n358), .A2(new_n365), .A3(new_n287), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT31), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  AND4_X1   g196(.A1(KEYINPUT31), .A2(new_n381), .A3(new_n378), .A4(new_n374), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n372), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n385));
  NOR2_X1   g199(.A1(G472), .A2(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT31), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n374), .A2(new_n378), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n381), .A2(KEYINPUT31), .A3(new_n378), .A4(new_n374), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n371), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n386), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT75), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G472), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n358), .A2(new_n365), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n378), .ZN(new_n400));
  INV_X1    g214(.A(new_n287), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n367), .A2(new_n370), .A3(new_n287), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n359), .A2(new_n375), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n358), .A2(new_n365), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n369), .B1(new_n407), .B2(KEYINPUT28), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n401), .A2(new_n404), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n266), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n398), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n393), .A2(new_n394), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(KEYINPUT32), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n280), .B1(new_n397), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(KEYINPUT71), .A2(G237), .ZN(new_n418));
  NOR2_X1   g232(.A1(KEYINPUT71), .A2(G237), .ZN(new_n419));
  OAI211_X1 g233(.A(G214), .B(new_n246), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n315), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n281), .A2(G143), .A3(G214), .A4(new_n246), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT88), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n421), .A2(new_n422), .A3(new_n427), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n421), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n421), .B2(new_n422), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n425), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n190), .B(new_n231), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n338), .B1(new_n421), .B2(new_n422), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n233), .B1(KEYINPUT17), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT17), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n422), .A3(new_n338), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n417), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n435), .A2(new_n442), .A3(new_n417), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT89), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n435), .A2(new_n442), .A3(new_n446), .A4(new_n417), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G475), .B1(new_n448), .B2(G902), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n438), .A2(new_n440), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n196), .B(KEYINPUT19), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n452), .B(new_n192), .C1(G146), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n435), .ZN(new_n455));
  INV_X1    g269(.A(new_n417), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n450), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n445), .A2(new_n447), .B1(new_n456), .B2(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(new_n459), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n461), .A2(KEYINPUT20), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n449), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT90), .B(new_n449), .C1(new_n460), .C2(new_n463), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n315), .A2(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n198), .A2(G143), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT93), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT93), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n331), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n294), .B2(G122), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT91), .A3(G116), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n295), .A2(G122), .A3(new_n296), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G107), .ZN(new_n483));
  INV_X1    g297(.A(G107), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n475), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n198), .A2(G143), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(KEYINPUT13), .B2(new_n469), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G134), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT92), .B1(new_n468), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT94), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n482), .B(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n490), .B(G134), .C1(new_n488), .C2(new_n493), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n475), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT95), .B1(new_n481), .B2(KEYINPUT14), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n480), .A3(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n481), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g319(.A(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n471), .A2(G134), .A3(new_n473), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n483), .B1(new_n475), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT9), .B(G234), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n510), .A2(new_n261), .A3(G953), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n501), .A2(KEYINPUT96), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n496), .A2(new_n500), .B1(new_n506), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT96), .B1(new_n513), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n262), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G478), .ZN(new_n517));
  NOR2_X1   g331(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(KEYINPUT97), .A2(KEYINPUT15), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n511), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n513), .ZN(new_n526));
  INV_X1    g340(.A(new_n511), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(new_n512), .ZN(new_n529));
  INV_X1    g343(.A(new_n521), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n262), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G952), .ZN(new_n533));
  AOI211_X1 g347(.A(G953), .B(new_n533), .C1(G234), .C2(G237), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n246), .B(new_n262), .C1(G234), .C2(G237), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n466), .A2(new_n467), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G122), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n416), .A2(G107), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n484), .A2(KEYINPUT3), .A3(G104), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT3), .B1(new_n484), .B2(G104), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G101), .ZN(new_n546));
  INV_X1    g360(.A(G101), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(KEYINPUT4), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT4), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n550), .A3(G101), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n306), .B2(new_n312), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n484), .B2(G104), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n484), .A2(G104), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n416), .A2(KEYINPUT83), .A3(G107), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G101), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n548), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n297), .A2(KEYINPUT5), .A3(new_n298), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(G113), .C1(KEYINPUT5), .C2(new_n298), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n311), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n541), .B1(new_n553), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n552), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT68), .B1(new_n311), .B2(new_n300), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n305), .B(new_n299), .C1(new_n309), .C2(new_n310), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n563), .A3(new_n540), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT6), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT6), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n541), .C1(new_n553), .C2(new_n564), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n324), .A2(new_n328), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G125), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(G125), .B2(new_n347), .ZN(new_n576));
  INV_X1    g390(.A(G224), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G953), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n576), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT7), .B1(new_n577), .B2(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n576), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n540), .B(KEYINPUT8), .Z(new_n583));
  NAND2_X1  g397(.A1(new_n311), .A2(new_n562), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n559), .A2(new_n548), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n586), .B2(new_n563), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n588), .B2(new_n570), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n580), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n580), .B2(new_n589), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G214), .B1(G237), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G221), .B1(new_n510), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G469), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n246), .A2(G227), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n560), .A2(KEYINPUT10), .A3(new_n347), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n317), .A2(new_n323), .A3(new_n319), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n343), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n585), .B1(new_n346), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n604), .B1(new_n607), .B2(KEYINPUT10), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n549), .A2(new_n329), .A3(new_n551), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n340), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT85), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n609), .B(new_n604), .C1(KEYINPUT10), .C2(new_n607), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n340), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n606), .A2(new_n346), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n585), .ZN(new_n619));
  INV_X1    g433(.A(new_n340), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n609), .A4(new_n604), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n603), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n560), .A2(new_n347), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n340), .B1(new_n623), .B2(new_n607), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT12), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n360), .A2(new_n585), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n618), .B2(new_n585), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n630), .A2(KEYINPUT84), .A3(new_n625), .A4(new_n340), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n621), .A2(new_n628), .A3(new_n631), .A4(new_n603), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n599), .B(new_n262), .C1(new_n622), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G902), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n599), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n614), .A2(new_n340), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n602), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n628), .A2(new_n631), .A3(new_n621), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n616), .A2(new_n637), .B1(new_n602), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n639), .B2(G469), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n598), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n596), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n539), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n414), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n526), .B2(new_n527), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n529), .A2(new_n646), .B1(new_n523), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n266), .A2(new_n517), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n648), .A2(new_n649), .B1(new_n517), .B2(new_n516), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n467), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT20), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n458), .A2(new_n653), .A3(new_n459), .ZN(new_n654));
  INV_X1    g468(.A(new_n450), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n461), .B2(new_n462), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT90), .B1(new_n657), .B2(new_n449), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n651), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n580), .A2(new_n589), .ZN(new_n660));
  INV_X1    g474(.A(new_n590), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n580), .A2(new_n589), .A3(new_n590), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n537), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n595), .B1(new_n592), .B2(KEYINPUT98), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n393), .B2(new_n266), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n387), .A2(new_n395), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n641), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n280), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT34), .B(G104), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  NAND3_X1  g491(.A1(new_n458), .A2(new_n459), .A3(new_n450), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n656), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n532), .A2(new_n679), .A3(new_n449), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n668), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n672), .A2(new_n674), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  INV_X1    g498(.A(new_n275), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT25), .B1(new_n259), .B2(new_n267), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n278), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n257), .A2(KEYINPUT36), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n256), .A2(KEYINPUT99), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n256), .A2(KEYINPUT99), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n688), .A3(new_n690), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n264), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n687), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n693), .A2(new_n695), .A3(new_n264), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT100), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n643), .A2(new_n672), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  NAND2_X1  g521(.A1(new_n397), .A2(new_n413), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n641), .A2(new_n665), .A3(new_n667), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(G900), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n534), .B1(new_n535), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n678), .B2(new_n656), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n449), .A3(new_n532), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n708), .A2(new_n704), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XNOR2_X1  g531(.A(new_n593), .B(KEYINPUT38), .ZN(new_n718));
  INV_X1    g532(.A(new_n532), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n687), .A2(new_n697), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n595), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n407), .A2(new_n401), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n389), .B2(new_n390), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n398), .B1(new_n723), .B2(new_n634), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n412), .B2(KEYINPUT32), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n397), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n712), .B(KEYINPUT39), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n641), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(KEYINPUT40), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n652), .A2(new_n658), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(KEYINPUT40), .B2(new_n728), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n721), .A2(new_n726), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  AOI211_X1 g547(.A(new_n650), .B(new_n712), .C1(new_n466), .C2(new_n467), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n708), .A2(new_n734), .A3(new_n704), .A4(new_n710), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  INV_X1    g550(.A(new_n632), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n636), .B1(new_n613), .B2(new_n615), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n603), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n599), .A2(KEYINPUT101), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n262), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n615), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT85), .B1(new_n614), .B2(new_n340), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n621), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n632), .B1(new_n745), .B2(new_n602), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n740), .B1(new_n746), .B2(new_n266), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n742), .A2(new_n747), .A3(new_n597), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n279), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n397), .B2(new_n413), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n669), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  INV_X1    g567(.A(new_n749), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n708), .A2(new_n681), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT102), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n757), .A3(new_n681), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  NAND3_X1  g574(.A1(new_n748), .A2(new_n665), .A3(new_n667), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n539), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n708), .A3(new_n704), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  OR2_X1    g578(.A1(new_n408), .A2(new_n287), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n382), .B2(new_n383), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n386), .B(KEYINPUT103), .Z(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n670), .A2(new_n768), .A3(new_n279), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n670), .A2(new_n768), .A3(new_n279), .A4(KEYINPUT104), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n665), .A2(new_n667), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n719), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n466), .A2(new_n467), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n742), .A2(new_n747), .A3(new_n597), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n537), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NAND3_X1  g595(.A1(new_n720), .A2(new_n670), .A3(new_n768), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n761), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n734), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n279), .A2(new_n641), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n708), .A2(new_n734), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT42), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n788), .B1(new_n397), .B2(new_n413), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n786), .B1(new_n793), .B2(new_n734), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n413), .B1(KEYINPUT32), .B2(new_n412), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n279), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n787), .A2(new_n641), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n797), .ZN(new_n798));
  OAI22_X1  g612(.A1(new_n792), .A2(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G131), .ZN(G33));
  AND2_X1   g614(.A1(new_n793), .A2(new_n715), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT106), .B(G134), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G36));
  NAND2_X1  g617(.A1(new_n730), .A2(new_n651), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT43), .Z(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n671), .A3(new_n720), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n639), .A2(KEYINPUT45), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n639), .A2(KEYINPUT45), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(G469), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT107), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n635), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n633), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(new_n597), .A3(new_n727), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n808), .A2(new_n787), .A3(new_n809), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n597), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(KEYINPUT47), .A3(new_n597), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n787), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n708), .A2(new_n279), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n734), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT108), .B(G140), .Z(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G42));
  NOR3_X1   g644(.A1(new_n720), .A2(new_n673), .A3(new_n712), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n726), .A2(new_n831), .A3(new_n776), .A4(new_n775), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n735), .A2(new_n716), .A3(new_n832), .A4(new_n784), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n703), .A2(new_n709), .A3(new_n714), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n835), .A2(new_n708), .B1(new_n783), .B2(new_n734), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n735), .A4(new_n832), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n466), .A2(new_n467), .A3(new_n532), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n659), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n596), .A2(new_n666), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n672), .A3(new_n674), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n846), .A2(new_n644), .A3(new_n705), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n797), .A2(new_n670), .A3(new_n720), .A4(new_n768), .ZN(new_n849));
  INV_X1    g663(.A(new_n712), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n776), .A2(new_n651), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n782), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n734), .A2(new_n853), .A3(KEYINPUT110), .A4(new_n797), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n522), .A2(new_n449), .A3(new_n531), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n787), .A2(new_n641), .A3(new_n713), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n703), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n715), .A2(new_n793), .B1(new_n858), .B2(new_n708), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n855), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n798), .A2(new_n796), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n790), .A2(new_n791), .ZN(new_n862));
  INV_X1    g676(.A(new_n794), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n757), .A2(new_n708), .A3(new_n681), .A4(new_n754), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n757), .B1(new_n750), .B2(new_n681), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n780), .A2(new_n751), .A3(new_n763), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n703), .A2(new_n761), .A3(new_n539), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n872), .A2(new_n708), .B1(new_n750), .B2(new_n669), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n780), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n834), .A2(KEYINPUT111), .A3(new_n838), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n841), .A2(new_n865), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n703), .A2(new_n671), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n643), .B1(new_n879), .B2(new_n414), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n846), .A2(new_n855), .A3(new_n880), .A4(new_n859), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n869), .A2(new_n870), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n799), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n878), .B1(new_n883), .B2(new_n839), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n841), .A2(new_n876), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT53), .B1(new_n883), .B2(new_n839), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n891), .B2(KEYINPUT54), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n805), .A2(new_n534), .A3(new_n773), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n595), .A3(new_n718), .A4(new_n748), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT50), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT50), .ZN(new_n898));
  INV_X1    g712(.A(new_n534), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n826), .A2(new_n777), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n805), .A2(new_n853), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n726), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n749), .A2(new_n899), .A3(new_n826), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n730), .A2(new_n650), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n742), .A2(new_n747), .A3(new_n598), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n823), .A2(new_n824), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n893), .A2(new_n787), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n897), .A2(new_n898), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n906), .B(KEYINPUT114), .Z(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n912), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n908), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n916), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n909), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n915), .A2(new_n919), .A3(new_n898), .A4(new_n897), .ZN(new_n920));
  INV_X1    g734(.A(new_n761), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n893), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT116), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n279), .A2(new_n805), .A3(new_n795), .A4(new_n900), .ZN(new_n924));
  AND2_X1   g738(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(G952), .B(new_n246), .C1(new_n904), .C2(new_n659), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n923), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n892), .A2(new_n913), .A3(new_n920), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(G952), .B2(G953), .ZN(new_n932));
  INV_X1    g746(.A(new_n718), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n742), .A2(new_n747), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT49), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n804), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n279), .A2(new_n597), .A3(new_n594), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n902), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n932), .A2(new_n939), .ZN(G75));
  NOR2_X1   g754(.A1(new_n246), .A2(G952), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n262), .B1(new_n877), .B2(new_n884), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT56), .B1(new_n943), .B2(new_n661), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n571), .A2(new_n573), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n579), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT55), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n942), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n944), .B2(new_n947), .ZN(G51));
  XNOR2_X1  g763(.A(new_n635), .B(KEYINPUT57), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n885), .B2(KEYINPUT54), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT54), .ZN(new_n953));
  AOI211_X1 g767(.A(KEYINPUT119), .B(new_n953), .C1(new_n877), .C2(new_n884), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT118), .B1(new_n885), .B2(KEYINPUT54), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n877), .A2(new_n884), .A3(new_n957), .A4(new_n953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT120), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n950), .C1(new_n955), .C2(new_n959), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n739), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n813), .B(KEYINPUT121), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n943), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n941), .B1(new_n964), .B2(new_n966), .ZN(G54));
  AND3_X1   g781(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n942), .B1(new_n968), .B2(new_n458), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n458), .B2(new_n968), .ZN(G60));
  INV_X1    g784(.A(new_n648), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n517), .A2(new_n634), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n892), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n648), .B(new_n974), .C1(new_n955), .C2(new_n959), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n942), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n877), .B2(new_n884), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n259), .A2(new_n260), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n942), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n696), .B2(new_n981), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n536), .B2(new_n577), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n882), .A2(new_n847), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n945), .B1(G898), .B2(new_n246), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  AOI21_X1  g804(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n728), .A2(new_n826), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n414), .A2(new_n843), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT124), .Z(new_n994));
  NAND3_X1  g808(.A1(new_n828), .A2(new_n819), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n836), .A2(new_n735), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n732), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT123), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n376), .A2(new_n377), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(new_n453), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1001), .A2(G953), .A3(new_n1003), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n796), .A2(new_n730), .A3(new_n719), .A4(new_n774), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n801), .B1(new_n818), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n828), .A2(new_n1006), .A3(new_n799), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n819), .A2(new_n996), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n819), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n246), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G900), .A2(G953), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n991), .B(new_n1004), .C1(new_n1015), .C2(new_n1003), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G227), .A2(G900), .ZN(new_n1017));
  AND4_X1   g831(.A1(G953), .A2(new_n1015), .A3(new_n1017), .A4(new_n1003), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1016), .A2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  OAI21_X1  g835(.A(new_n402), .B1(new_n389), .B2(new_n390), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n891), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1021), .B(KEYINPUT126), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n1001), .B2(new_n987), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n400), .A2(new_n287), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1025), .B1(new_n1012), .B2(new_n987), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n399), .A2(new_n401), .A3(new_n378), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n942), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(KEYINPUT127), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1033), .B(new_n942), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1028), .B1(new_n1032), .B2(new_n1034), .ZN(G57));
endmodule


