//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT90), .B(G224), .Z(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT7), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT0), .B(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT72), .A2(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n195), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n193), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G128), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT92), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g029(.A(KEYINPUT92), .B(new_n205), .C1(new_n210), .C2(new_n212), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n192), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT93), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT93), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(new_n192), .C1(new_n215), .C2(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n224), .A3(G104), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n228), .A2(new_n224), .A3(KEYINPUT3), .A4(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G101), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n224), .B2(G104), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(KEYINPUT82), .A3(new_n236), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n227), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  OAI21_X1  g057(.A(G113), .B1(new_n243), .B2(KEYINPUT5), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n242), .A2(G116), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT67), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(G119), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n243), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n244), .B1(new_n252), .B2(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(new_n249), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n241), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT81), .B1(new_n263), .B2(new_n234), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT82), .B1(new_n233), .B2(new_n236), .ZN(new_n265));
  AOI211_X1 g079(.A(new_n238), .B(new_n235), .C1(new_n231), .C2(new_n232), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT3), .B1(new_n223), .B2(new_n228), .ZN(new_n268));
  INV_X1    g082(.A(new_n232), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n268), .A2(new_n269), .B1(G104), .B2(new_n224), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G101), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT4), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n248), .A2(new_n255), .A3(new_n251), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n256), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT68), .B1(new_n275), .B2(new_n256), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n270), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n263), .A2(KEYINPUT83), .A3(new_n281), .ZN(new_n282));
  OAI22_X1  g096(.A1(new_n276), .A2(new_n277), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n259), .B(new_n262), .C1(new_n274), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n213), .B1(new_n206), .B2(KEYINPUT89), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(KEYINPUT89), .B2(new_n206), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n286), .A2(new_n192), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n221), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n226), .B1(new_n265), .B2(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n258), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n239), .A2(new_n240), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n243), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n256), .B1(new_n292), .B2(new_n244), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n226), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n262), .B(KEYINPUT8), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT91), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n288), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n259), .B1(new_n274), .B2(new_n283), .ZN(new_n300));
  INV_X1    g114(.A(new_n262), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n286), .B(new_n191), .Z(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT94), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n299), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n299), .B2(new_n307), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n190), .A2(G952), .ZN(new_n316));
  NAND2_X1  g130(.A1(G234), .A2(G237), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(G902), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT21), .B(G898), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n313), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n190), .A2(G227), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n326), .B(new_n327), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n272), .A4(new_n264), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n270), .A2(new_n278), .A3(new_n279), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT83), .B1(new_n263), .B2(new_n281), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n200), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n210), .A2(new_n212), .A3(new_n226), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n265), .B2(new_n266), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT10), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n334), .C1(new_n265), .C2(new_n266), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n330), .A2(new_n333), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G134), .ZN(new_n341));
  INV_X1    g155(.A(G134), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT11), .B1(new_n342), .B2(G137), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n340), .A3(G134), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n341), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G131), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(KEYINPUT64), .A3(new_n347), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT84), .B1(new_n339), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n336), .A2(new_n338), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n333), .B1(new_n267), .B2(new_n273), .ZN(new_n358));
  AND4_X1   g172(.A1(KEYINPUT84), .A2(new_n357), .A3(new_n358), .A4(new_n355), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n329), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT12), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n210), .A2(new_n212), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(new_n289), .B1(new_n291), .B2(new_n334), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  INV_X1    g178(.A(new_n362), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n335), .B1(new_n241), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n346), .A2(new_n347), .ZN(new_n367));
  AND4_X1   g181(.A1(KEYINPUT64), .A2(new_n349), .A3(new_n347), .A4(new_n350), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT64), .B1(new_n346), .B2(new_n347), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(KEYINPUT85), .A3(KEYINPUT12), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n289), .A2(new_n362), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n355), .B1(new_n373), .B2(new_n335), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT85), .B1(new_n374), .B2(KEYINPUT12), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n325), .B1(new_n360), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n357), .A2(new_n358), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n370), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n339), .A2(KEYINPUT84), .A3(new_n355), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n366), .A2(KEYINPUT12), .A3(new_n370), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n364), .A3(new_n371), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT87), .A4(new_n329), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n356), .B2(new_n359), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n328), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n377), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  INV_X1    g207(.A(G902), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n329), .B1(new_n382), .B2(new_n386), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n328), .B(new_n388), .C1(new_n380), .C2(new_n381), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT86), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n382), .A2(new_n329), .A3(new_n389), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n364), .A2(new_n371), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n401), .A2(new_n385), .B1(new_n380), .B2(new_n381), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n399), .B(new_n400), .C1(new_n402), .C2(new_n329), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n403), .A3(G469), .ZN(new_n404));
  NAND2_X1  g218(.A1(G469), .A2(G902), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n395), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G217), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n187), .A2(new_n407), .A3(G953), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT100), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT97), .B1(new_n195), .B2(G128), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT97), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n211), .A3(G143), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n195), .A2(G128), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n413), .A2(KEYINPUT99), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT99), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n342), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G116), .B(G122), .Z(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(G107), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT13), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n410), .A2(new_n412), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(KEYINPUT98), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n414), .A2(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n422), .B2(KEYINPUT98), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n342), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n409), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n414), .A2(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n413), .A2(KEYINPUT98), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n421), .B2(new_n414), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n422), .A2(KEYINPUT98), .ZN(new_n431));
  OAI21_X1  g245(.A(G134), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT100), .A3(new_n417), .A4(new_n419), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n245), .A2(G122), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n224), .B1(new_n435), .B2(KEYINPUT14), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(new_n418), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n413), .A2(new_n414), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT99), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n413), .A2(KEYINPUT99), .A3(new_n414), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(G134), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n437), .B1(new_n417), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n408), .B1(new_n434), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n408), .ZN(new_n446));
  AOI211_X1 g260(.A(new_n443), .B(new_n446), .C1(new_n427), .C2(new_n433), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n394), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G478), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n449), .A2(KEYINPUT15), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n448), .B(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT96), .B(G475), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n203), .A2(G140), .A3(new_n204), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT71), .B1(new_n202), .B2(G140), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n456));
  INV_X1    g270(.A(G140), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G125), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(KEYINPUT16), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT73), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n455), .A2(new_n458), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT16), .A4(new_n454), .ZN(new_n463));
  NOR2_X1   g277(.A1(KEYINPUT16), .A2(G140), .ZN(new_n464));
  INV_X1    g278(.A(new_n204), .ZN(new_n465));
  NOR2_X1   g279(.A1(KEYINPUT72), .A2(G125), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT74), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT74), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n205), .A2(new_n469), .A3(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n193), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n460), .A2(new_n471), .A3(new_n463), .A4(G146), .ZN(new_n474));
  NOR2_X1   g288(.A1(G237), .A2(G953), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n475), .A2(G143), .A3(G214), .ZN(new_n476));
  AOI21_X1  g290(.A(G143), .B1(new_n475), .B2(G214), .ZN(new_n477));
  OAI21_X1  g291(.A(G131), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n479));
  INV_X1    g293(.A(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n190), .A3(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n195), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(G143), .A3(G214), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n347), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT17), .A3(G131), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n473), .A2(new_n474), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n486), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n457), .A2(G125), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n202), .A2(G140), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT77), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n492), .B2(new_n493), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G146), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n193), .B1(new_n461), .B2(new_n454), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G113), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(new_n222), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n503), .A3(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n453), .B1(new_n507), .B2(new_n394), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n489), .A2(new_n503), .A3(new_n500), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n461), .A2(new_n454), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT19), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n495), .B2(new_n496), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n193), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n474), .A2(new_n514), .A3(KEYINPUT95), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n478), .A2(new_n484), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT95), .B1(new_n474), .B2(new_n514), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n500), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n509), .B1(new_n504), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  INV_X1    g338(.A(new_n518), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n516), .A3(new_n515), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n503), .B1(new_n526), .B2(new_n500), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n524), .B(new_n521), .C1(new_n527), .C2(new_n509), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n508), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n451), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AND4_X1   g345(.A1(new_n188), .A2(new_n324), .A3(new_n406), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n368), .A2(new_n369), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n350), .A2(KEYINPUT66), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n342), .A3(G137), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT65), .B1(new_n342), .B2(G137), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT65), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n340), .A3(G134), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G131), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n212), .A3(new_n210), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n355), .A2(new_n200), .B1(new_n533), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n277), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n256), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n200), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n370), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n362), .B1(G131), .B2(new_n540), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n353), .A2(new_n354), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n549), .A2(new_n552), .B1(new_n544), .B2(new_n545), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT28), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n475), .A2(G210), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT27), .Z(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT26), .B(G101), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n276), .A2(new_n277), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n549), .A2(new_n560), .A3(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n543), .A2(KEYINPUT30), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT30), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n567), .A3(new_n552), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n547), .B1(new_n569), .B2(new_n546), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n564), .B(new_n565), .C1(new_n570), .C2(new_n559), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(new_n394), .C1(new_n565), .C2(new_n564), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n546), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n561), .A3(new_n559), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT31), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n543), .A2(new_n546), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n562), .B1(new_n577), .B2(new_n561), .ZN(new_n578));
  INV_X1    g392(.A(new_n543), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT28), .B1(new_n579), .B2(new_n560), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n558), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT69), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n583), .A3(new_n559), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n558), .C1(new_n578), .C2(new_n580), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n576), .A2(new_n582), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NOR2_X1   g402(.A1(G472), .A2(G902), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n573), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT23), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n242), .B2(G128), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n594), .B(new_n595), .C1(G119), .C2(new_n211), .ZN(new_n596));
  OR3_X1    g410(.A1(new_n596), .A2(KEYINPUT76), .A3(G110), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT76), .B1(new_n596), .B2(G110), .ZN(new_n598));
  XOR2_X1   g412(.A(G119), .B(G128), .Z(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT24), .B(G110), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n597), .B(new_n598), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n603), .B(new_n474), .C1(G146), .C2(new_n497), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n473), .A2(new_n474), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n600), .A2(new_n602), .B1(new_n596), .B2(G110), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT75), .B(new_n609), .C1(new_n473), .C2(new_n474), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n604), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT78), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(KEYINPUT78), .B(new_n604), .C1(new_n608), .C2(new_n610), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT79), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT22), .B(G137), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n604), .B(new_n618), .C1(new_n608), .C2(new_n610), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G234), .ZN(new_n623));
  OAI21_X1  g437(.A(G217), .B1(new_n623), .B2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n394), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n624), .B(KEYINPUT70), .Z(new_n627));
  AND2_X1   g441(.A1(new_n621), .A2(new_n394), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n629), .B2(KEYINPUT25), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT25), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n620), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n626), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n592), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n532), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  INV_X1    g451(.A(new_n633), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n587), .B2(new_n394), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n587), .A2(new_n589), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n640), .B2(KEYINPUT101), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n406), .A2(new_n188), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n299), .A2(new_n307), .A3(KEYINPUT102), .A4(new_n310), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n314), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n313), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n323), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n434), .A2(new_n444), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n446), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n434), .A2(new_n444), .A3(new_n408), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT33), .B1(new_n445), .B2(new_n447), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(G478), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n449), .B(new_n394), .C1(new_n445), .C2(new_n447), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n449), .A2(new_n394), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n529), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n650), .A2(new_n651), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n644), .A2(new_n646), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT103), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND2_X1  g482(.A1(new_n523), .A2(new_n528), .ZN(new_n669));
  INV_X1    g483(.A(new_n508), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n451), .ZN(new_n672));
  INV_X1    g486(.A(new_n648), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n296), .B(KEYINPUT91), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n221), .A2(new_n284), .A3(new_n287), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n394), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n309), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n299), .A2(new_n307), .A3(new_n310), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n649), .A3(new_n679), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n651), .A2(new_n672), .A3(new_n673), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n644), .A2(new_n646), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  OR2_X1    g498(.A1(new_n619), .A2(KEYINPUT36), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n613), .A2(new_n614), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n613), .B2(new_n614), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n625), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n630), .B2(new_n632), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n641), .A2(new_n643), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n532), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT37), .B(G110), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT104), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n691), .B(new_n693), .ZN(G12));
  NAND2_X1  g508(.A1(new_n629), .A2(KEYINPUT25), .ZN(new_n695));
  INV_X1    g509(.A(new_n627), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n632), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n688), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n592), .A2(new_n650), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n451), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n320), .A2(G900), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n318), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n529), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n700), .A2(new_n646), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n703), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n646), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n570), .A2(new_n558), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n577), .A2(new_n561), .A3(new_n558), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n394), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n590), .B2(new_n591), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n689), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n313), .B(new_n717), .Z(new_n718));
  NOR2_X1   g532(.A1(new_n451), .A2(new_n529), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n314), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n710), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n663), .B2(new_n703), .ZN(new_n725));
  INV_X1    g539(.A(new_n703), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n662), .A2(new_n529), .A3(KEYINPUT106), .A4(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n700), .A2(new_n646), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  NAND2_X1  g544(.A1(new_n392), .A2(new_n394), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n188), .A3(new_n395), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n634), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n664), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT107), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n736), .B(new_n738), .ZN(G15));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n681), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  AND4_X1   g555(.A1(new_n188), .A2(new_n650), .A3(new_n395), .A4(new_n732), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n530), .A2(new_n323), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n592), .A2(new_n699), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND3_X1  g560(.A1(new_n576), .A2(new_n584), .A3(new_n581), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n589), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n554), .A2(new_n563), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n585), .B1(new_n749), .B2(new_n558), .ZN(new_n750));
  INV_X1    g564(.A(new_n586), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n583), .B1(new_n570), .B2(new_n559), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n560), .B1(new_n566), .B2(new_n568), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n547), .A4(new_n558), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(G902), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n748), .B1(new_n757), .B2(new_n639), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n638), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n701), .A2(new_n760), .A3(new_n671), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n451), .B2(new_n529), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n680), .A2(new_n761), .A3(new_n762), .A4(new_n673), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n759), .A2(new_n763), .A3(new_n733), .A4(new_n651), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NOR2_X1   g579(.A1(new_n689), .A2(new_n758), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n728), .A2(new_n733), .A3(new_n650), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  INV_X1    g583(.A(new_n188), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n315), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n678), .A2(new_n679), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n396), .A2(new_n397), .ZN(new_n773));
  OAI21_X1  g587(.A(G469), .B1(new_n773), .B2(G902), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n395), .B2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n775), .A2(new_n592), .A3(new_n633), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n659), .A2(new_n661), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n671), .A2(new_n658), .A3(new_n778), .A4(new_n703), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT106), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n663), .A2(new_n724), .A3(new_n703), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n769), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n728), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT109), .B(G131), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G33));
  XNOR2_X1  g601(.A(new_n704), .B(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n776), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND2_X1  g604(.A1(new_n773), .A2(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(G469), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n398), .B2(new_n403), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n405), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n395), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n770), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n708), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n529), .A2(new_n658), .A3(new_n778), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT43), .Z(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(new_n699), .C1(new_n641), .C2(new_n643), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n800), .B(new_n807), .C1(new_n806), .C2(new_n805), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  NOR4_X1   g623(.A1(new_n782), .A2(new_n633), .A3(new_n592), .A4(new_n802), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NOR4_X1   g628(.A1(new_n718), .A2(new_n770), .A3(new_n315), .A4(new_n803), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n638), .A2(new_n715), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n732), .A2(new_n395), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT49), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n678), .A2(new_n679), .A3(new_n314), .A4(new_n703), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n530), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n592), .A2(new_n821), .A3(new_n699), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n776), .A2(new_n788), .B1(new_n822), .B2(new_n646), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n395), .A2(new_n774), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n747), .A2(new_n589), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n640), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n772), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n699), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT114), .B1(new_n828), .B2(new_n782), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n728), .A2(new_n830), .A3(new_n766), .A4(new_n775), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n823), .A2(new_n832), .A3(KEYINPUT115), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(new_n836), .B1(new_n783), .B2(new_n784), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n592), .A2(new_n650), .A3(new_n699), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n645), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n699), .A2(new_n826), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n782), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n839), .A2(new_n705), .B1(new_n841), .B2(new_n742), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n703), .B(KEYINPUT116), .Z(new_n844));
  AND4_X1   g658(.A1(new_n697), .A2(new_n698), .A3(new_n188), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n763), .A2(new_n845), .A3(new_n715), .A4(new_n824), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(new_n843), .A3(new_n729), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n706), .A2(new_n729), .A3(new_n767), .A4(new_n846), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n671), .B2(new_n451), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n671), .A2(new_n451), .A3(KEYINPUT112), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n324), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n324), .A2(new_n855), .A3(new_n851), .A4(new_n852), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n644), .A3(new_n646), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n532), .B1(new_n635), .B2(new_n690), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n644), .A2(new_n646), .A3(new_n324), .A4(new_n663), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n635), .B(new_n733), .C1(new_n664), .C2(new_n681), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n745), .A3(new_n764), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(new_n745), .A3(new_n764), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n837), .A2(new_n850), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n843), .B1(new_n706), .B2(new_n767), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT53), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n823), .A2(new_n832), .A3(KEYINPUT115), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT115), .B1(new_n823), .B2(new_n832), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n785), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n847), .A2(new_n849), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n875), .B2(new_n866), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n861), .A2(new_n745), .A3(new_n764), .A4(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n860), .A2(new_n881), .A3(new_n868), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n837), .A2(new_n850), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n817), .A2(new_n319), .A3(new_n827), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n816), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n529), .A3(new_n662), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n804), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n840), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n734), .A2(new_n718), .A3(new_n314), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n759), .A2(new_n804), .A3(new_n319), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT50), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(KEYINPUT50), .A3(new_n892), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n812), .B(new_n811), .C1(new_n770), .C2(new_n817), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n801), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(new_n887), .ZN(new_n903));
  INV_X1    g717(.A(new_n663), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n316), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n889), .A2(new_n634), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT48), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n905), .B(new_n907), .C1(new_n742), .C2(new_n892), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n885), .A2(new_n901), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n819), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n190), .A2(G952), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT118), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n394), .B1(new_n879), .B2(new_n883), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(new_n309), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n303), .A2(new_n305), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT117), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n306), .B(KEYINPUT55), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(new_n921));
  OR2_X1    g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n921), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(G51));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n883), .A2(new_n880), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n876), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n883), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n876), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n879), .A2(KEYINPUT120), .A3(new_n880), .A4(new_n883), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n405), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n392), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n792), .A2(new_n793), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n916), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n913), .B1(new_n935), .B2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(new_n520), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n520), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n913), .ZN(G60));
  NAND2_X1  g756(.A1(new_n656), .A2(new_n657), .ZN(new_n943));
  XNOR2_X1  g757(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n661), .B(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n931), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n877), .B2(new_n884), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n914), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n879), .B2(new_n883), .ZN(new_n953));
  INV_X1    g767(.A(new_n622), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n686), .A2(new_n687), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n914), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(new_n189), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n963), .B2(new_n322), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n866), .B2(G953), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n919), .B1(G898), .B2(new_n190), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT122), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  AOI21_X1  g782(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n511), .A2(new_n513), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n569), .B(new_n970), .Z(new_n971));
  NAND3_X1  g785(.A1(new_n722), .A2(new_n729), .A3(new_n842), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n975), .A3(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n808), .A2(new_n813), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n722), .A2(new_n979), .A3(new_n729), .A4(new_n842), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n635), .A2(new_n801), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n852), .A2(new_n851), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n709), .B(new_n981), .C1(new_n904), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n977), .A2(new_n978), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n971), .B1(new_n986), .B2(new_n190), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n635), .A2(new_n763), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n800), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT126), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n729), .A2(new_n785), .A3(new_n789), .A4(new_n842), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n978), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(G900), .A2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n971), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n969), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n993), .A2(new_n995), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n969), .B(KEYINPUT125), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT124), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n998), .B(new_n999), .C1(new_n987), .C2(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n987), .A2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  NAND2_X1  g819(.A1(new_n863), .A2(new_n865), .ZN(new_n1006));
  INV_X1    g820(.A(new_n860), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1005), .B1(new_n992), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n570), .A2(new_n558), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n913), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1005), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n985), .A2(new_n978), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n976), .B2(new_n974), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1013), .B1(new_n1015), .B2(new_n866), .ZN(new_n1016));
  INV_X1    g830(.A(new_n711), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n870), .A2(new_n876), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n1010), .A3(new_n1005), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(G57));
endmodule


