//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n208), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT73), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(KEYINPUT73), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n202), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT3), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G155gat), .B(G162gat), .Z(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n224), .A2(new_n229), .A3(KEYINPUT2), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(new_n221), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n223), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(KEYINPUT78), .A3(new_n223), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n218), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  INV_X1    g039(.A(new_n227), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n231), .A2(KEYINPUT78), .A3(new_n223), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT78), .B1(new_n231), .B2(new_n223), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n217), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n207), .B1(new_n206), .B2(new_n208), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n202), .B1(new_n246), .B2(new_n214), .ZN(new_n247));
  INV_X1    g046(.A(new_n215), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT74), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT74), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n213), .A2(new_n250), .A3(new_n215), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT81), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT31), .B(G50gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n239), .A2(new_n253), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n218), .B2(new_n236), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n213), .B2(new_n215), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n262), .B(KEYINPUT82), .C1(new_n263), .C2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n253), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n265), .A2(new_n266), .A3(new_n238), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n265), .B2(new_n238), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n258), .A2(new_n254), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT85), .B(G22gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n270), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n273), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n271), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n278), .A2(KEYINPUT23), .B1(new_n281), .B2(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G183gat), .B(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n290), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT25), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G190gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT24), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(KEYINPUT23), .B2(new_n278), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n301), .A2(new_n291), .A3(new_n303), .A4(new_n294), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n305));
  AOI22_X1  g104(.A1(new_n289), .A2(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n281), .ZN(new_n310));
  NOR3_X1   g109(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n307), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(new_n297), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(new_n297), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n312), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n278), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(new_n281), .A3(new_n309), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n307), .B1(new_n324), .B2(new_n308), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G226gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n306), .A2(new_n326), .B1(KEYINPUT29), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n304), .A2(new_n305), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n287), .B1(new_n286), .B2(new_n280), .ZN(new_n332));
  AND4_X1   g131(.A1(new_n287), .A2(new_n279), .A3(new_n280), .A4(new_n283), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n291), .A4(new_n294), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n325), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(new_n312), .A3(new_n315), .A4(new_n320), .ZN(new_n338));
  INV_X1    g137(.A(new_n329), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n252), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n249), .A2(new_n251), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n330), .A3(new_n340), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT30), .A4(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT76), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n343), .A2(new_n330), .A3(new_n340), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n330), .A2(new_n340), .B1(new_n249), .B2(new_n251), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n342), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n347), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n357), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n349), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G227gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n328), .ZN(new_n364));
  XNOR2_X1  g163(.A(G127gat), .B(G134gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G113gat), .A2(G120gat), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n365), .A2(new_n366), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(G113gat), .A2(G120gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT69), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n376), .A3(new_n370), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n377), .A3(new_n366), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT68), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G127gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n365), .A2(new_n379), .B1(G134gat), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT70), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n372), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n306), .B2(new_n326), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n378), .A2(new_n381), .A3(new_n384), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n378), .B2(new_n381), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n371), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n336), .A3(new_n338), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n364), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI211_X1 g193(.A(KEYINPUT34), .B(new_n364), .C1(new_n387), .C2(new_n391), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n364), .A3(new_n391), .ZN(new_n397));
  XOR2_X1   g196(.A(G71gat), .B(G99gat), .Z(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT33), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT71), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(KEYINPUT32), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n387), .A2(new_n391), .A3(new_n364), .A4(new_n400), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n406), .B2(new_n401), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n396), .B(new_n404), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n405), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n394), .A2(new_n395), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT89), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n362), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT35), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n418));
  NAND2_X1  g217(.A1(new_n386), .A2(new_n236), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n390), .A2(new_n262), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n244), .A3(new_n390), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n390), .B2(new_n262), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n386), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n426), .A2(new_n422), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n390), .A2(new_n262), .A3(new_n427), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT4), .B1(new_n386), .B2(new_n236), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(new_n418), .A3(new_n422), .A4(new_n426), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n435), .A3(new_n440), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT86), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n440), .B(new_n443), .C1(new_n431), .C2(new_n435), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n431), .B2(new_n435), .ZN(new_n449));
  INV_X1    g248(.A(new_n443), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n444), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n277), .A2(new_n416), .A3(new_n417), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n272), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n265), .A2(new_n238), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n265), .A2(new_n266), .A3(new_n238), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n273), .B1(new_n460), .B2(new_n259), .ZN(new_n461));
  INV_X1    g260(.A(new_n274), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n404), .C1(new_n407), .C2(new_n405), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(new_n410), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n362), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n445), .A2(new_n448), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n423), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(KEYINPUT39), .C1(new_n423), .C2(new_n421), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n477), .A3(new_n423), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n440), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n449), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n362), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n464), .A3(new_n463), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n344), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n359), .B2(new_n485), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n342), .A2(new_n488), .A3(new_n344), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n357), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n487), .A2(new_n491), .B1(new_n360), .B2(new_n357), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n447), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n446), .A2(new_n453), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n356), .A2(KEYINPUT37), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n357), .A3(new_n489), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n494), .A2(new_n495), .B1(KEYINPUT38), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n446), .A2(new_n493), .A3(new_n453), .A4(KEYINPUT88), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n447), .B1(new_n451), .B2(new_n444), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n275), .A2(new_n276), .B1(new_n501), .B2(new_n362), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n467), .A2(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n408), .A2(new_n411), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n473), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G50gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(G43gat), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n514), .A2(new_n515), .A3(G50gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT15), .B1(new_n515), .B2(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n515), .B2(G50gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G29gat), .A2(G36gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT14), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n512), .A2(new_n520), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n522), .B1(new_n511), .B2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n532), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(G8gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(G8gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n531), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n537), .A2(KEYINPUT93), .A3(new_n538), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT93), .B1(new_n537), .B2(new_n538), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n529), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n547), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n545), .A2(new_n546), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n530), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n547), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n544), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT11), .B(G169gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT12), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n550), .A2(new_n556), .A3(new_n564), .A4(new_n551), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G231gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(new_n328), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569));
  INV_X1    g368(.A(G71gat), .ZN(new_n570));
  INV_X1    g369(.A(G78gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G78gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT96), .B(G57gat), .Z(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n575), .A2(G57gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n573), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n575), .A2(G57gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n572), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n580), .A2(KEYINPUT95), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT95), .B1(new_n580), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n568), .B1(new_n586), .B2(KEYINPUT21), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n585), .B(new_n588), .C1(new_n567), .C2(new_n328), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G127gat), .ZN(new_n591));
  INV_X1    g390(.A(G127gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n552), .B1(new_n588), .B2(new_n585), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  INV_X1    g398(.A(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n597), .B2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT7), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n531), .A2(new_n542), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n620), .A2(KEYINPUT97), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n529), .B2(new_n617), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(KEYINPUT97), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n621), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n585), .A2(new_n618), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n617), .B(new_n578), .C1(new_n583), .C2(new_n584), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n641), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n638), .B2(new_n639), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT98), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n641), .B1(new_n635), .B2(new_n637), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n644), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n646), .B2(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n608), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n508), .A2(new_n566), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n501), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(new_n362), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n362), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G8gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n663), .ZN(new_n666));
  MUX2_X1   g465(.A(new_n663), .B(new_n666), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT89), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT89), .B1(new_n408), .B2(new_n411), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n659), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n503), .A2(new_n505), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n676), .B2(new_n668), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n463), .A2(new_n464), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n659), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n566), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n607), .A2(new_n682), .A3(new_n656), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n508), .A2(new_n634), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n501), .A3(new_n509), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n683), .B(KEYINPUT99), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n494), .A2(new_n495), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n497), .A2(KEYINPUT38), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n499), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n484), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n507), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n463), .A2(new_n417), .A3(new_n464), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n469), .B1(new_n669), .B2(new_n670), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n501), .A2(new_n362), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(new_n464), .A3(new_n463), .A4(new_n467), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n696), .A2(new_n454), .B1(new_n698), .B2(KEYINPUT35), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n634), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n502), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n471), .A3(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n506), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n473), .B1(new_n705), .B2(new_n500), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n633), .A2(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n688), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n470), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n687), .B1(new_n509), .B2(new_n711), .ZN(G1328gat));
  NOR3_X1   g511(.A1(new_n684), .A2(G36gat), .A3(new_n469), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT46), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n710), .B2(new_n469), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n672), .A2(new_n515), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n684), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n683), .B(KEYINPUT99), .Z(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n508), .B2(new_n634), .ZN(new_n722));
  INV_X1    g521(.A(new_n707), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n691), .A2(new_n692), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n463), .A2(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n674), .B1(new_n725), .B2(KEYINPUT100), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(new_n703), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n723), .B1(new_n727), .B2(new_n473), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n674), .B(new_n720), .C1(new_n722), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n719), .B1(new_n729), .B2(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n717), .B1(new_n730), .B2(KEYINPUT47), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n515), .B1(new_n709), .B2(new_n674), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT101), .B(new_n732), .C1(new_n733), .C2(new_n719), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT47), .B1(new_n684), .B2(new_n718), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n515), .B1(new_n729), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n701), .A2(new_n708), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n740), .A2(KEYINPUT102), .A3(new_n674), .A4(new_n720), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n736), .B(new_n737), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n729), .A2(new_n738), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(G43gat), .A3(new_n741), .ZN(new_n744));
  INV_X1    g543(.A(new_n737), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT103), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n735), .B1(new_n742), .B2(new_n746), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n685), .B2(new_n678), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(KEYINPUT104), .B2(KEYINPUT48), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n709), .A2(G50gat), .A3(new_n678), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1331gat));
  NAND4_X1  g552(.A1(new_n607), .A2(new_n682), .A3(new_n633), .A4(new_n656), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n473), .B2(new_n727), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n501), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT105), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(new_n574), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n362), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  NAND3_X1  g561(.A1(new_n755), .A2(G71gat), .A3(new_n674), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n755), .A2(new_n672), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n765), .A2(new_n766), .B1(G71gat), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n755), .A2(new_n678), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n607), .A2(new_n566), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n706), .A2(new_n634), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n633), .B1(new_n727), .B2(new_n473), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(KEYINPUT108), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n772), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n773), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n774), .A2(new_n775), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n612), .A3(new_n501), .A4(new_n656), .ZN(new_n785));
  INV_X1    g584(.A(new_n656), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n786), .B(new_n780), .C1(new_n701), .C2(new_n708), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n501), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G85gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n469), .A2(new_n786), .A3(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n779), .B2(new_n783), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n613), .B1(new_n787), .B2(new_n362), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n796), .B2(new_n799), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1337gat));
  NOR3_X1   g602(.A1(new_n671), .A2(new_n786), .A3(G99gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n674), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1338gat));
  INV_X1    g607(.A(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n678), .A2(new_n809), .A3(new_n656), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT109), .Z(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n779), .B2(new_n783), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n809), .B1(new_n787), .B2(new_n678), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n813), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1339gat));
  NAND3_X1  g619(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n644), .A2(new_n822), .A3(new_n647), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n651), .B1(new_n646), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n825), .A3(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n654), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT110), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n829), .A3(new_n654), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n825), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n828), .A2(new_n566), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n554), .A2(new_n555), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n544), .B1(new_n543), .B2(new_n547), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n561), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n656), .A2(new_n565), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n634), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  AND4_X1   g638(.A1(new_n565), .A2(new_n631), .A3(new_n632), .A4(new_n837), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n828), .A3(new_n830), .A4(new_n833), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n608), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n607), .A2(new_n682), .A3(new_n633), .A4(new_n786), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n678), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n501), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n469), .A2(new_n467), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n367), .A3(new_n566), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n501), .A3(new_n416), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n845), .A2(KEYINPUT111), .A3(new_n501), .A4(new_n416), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n566), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n854), .A2(new_n855), .A3(G113gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n854), .B2(G113gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n848), .B2(new_n656), .ZN(new_n859));
  AND4_X1   g658(.A1(G120gat), .A2(new_n852), .A3(new_n656), .A4(new_n853), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n848), .A2(new_n592), .A3(new_n607), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n852), .A2(new_n607), .A3(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n592), .ZN(G1342gat));
  NOR2_X1   g663(.A1(new_n633), .A2(G134gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n847), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT56), .Z(new_n867));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n634), .A3(new_n853), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G134gat), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n674), .A2(new_n470), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n469), .ZN(new_n872));
  INV_X1    g671(.A(new_n831), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n874));
  OAI21_X1  g673(.A(new_n566), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n838), .B1(new_n875), .B2(new_n827), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n633), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n607), .B1(new_n877), .B2(new_n841), .ZN(new_n878));
  INV_X1    g677(.A(new_n844), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n678), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n872), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n843), .A2(new_n844), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n678), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n682), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n277), .B1(new_n843), .B2(new_n844), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n682), .A2(G141gat), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT114), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n889), .A2(new_n872), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n871), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT115), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(KEYINPUT115), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n362), .B(new_n891), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n897), .B2(new_n899), .ZN(G1344gat));
  XNOR2_X1  g699(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n901));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n883), .B(new_n678), .C1(new_n878), .C2(new_n879), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n872), .A2(new_n786), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n903), .B(new_n904), .C1(new_n888), .C2(new_n883), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n906), .B2(KEYINPUT119), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n901), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n881), .A2(new_n884), .A3(new_n656), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n902), .A2(KEYINPUT59), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n896), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n469), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n656), .A2(new_n902), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n910), .A2(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n885), .B2(new_n608), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n607), .A2(new_n600), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n918), .B2(new_n922), .ZN(G1346gat));
  NOR2_X1   g722(.A1(new_n885), .A2(new_n633), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT120), .ZN(new_n925));
  OAI21_X1  g724(.A(G162gat), .B1(new_n924), .B2(KEYINPUT120), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n633), .A2(G162gat), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n925), .A2(new_n926), .B1(new_n918), .B2(new_n927), .ZN(G1347gat));
  AOI21_X1  g727(.A(new_n501), .B1(new_n843), .B2(new_n844), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n468), .A2(new_n469), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n682), .A2(G169gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n470), .A2(new_n362), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT122), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n671), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n845), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n682), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n935), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n940), .B2(new_n786), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n932), .A2(new_n933), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n786), .A2(G176gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1349gat));
  NOR2_X1   g747(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n949));
  OAI21_X1  g748(.A(G183gat), .B1(new_n940), .B2(new_n608), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n929), .A2(new_n313), .A3(new_n607), .A4(new_n930), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n952), .B(new_n953), .Z(G1350gat));
  OAI21_X1  g753(.A(G190gat), .B1(new_n940), .B2(new_n633), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n634), .A2(new_n297), .ZN(new_n958));
  OAI22_X1  g757(.A1(new_n956), .A2(new_n957), .B1(new_n946), .B2(new_n958), .ZN(G1351gat));
  NAND3_X1  g758(.A1(new_n506), .A2(new_n678), .A3(new_n362), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n929), .A2(new_n961), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n962), .A2(G197gat), .A3(new_n682), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n938), .A2(new_n674), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n903), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n966), .B2(new_n682), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G197gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n966), .A2(KEYINPUT126), .A3(new_n682), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  NOR2_X1   g769(.A1(new_n786), .A2(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n962), .A2(KEYINPUT127), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(new_n962), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G204gat), .B1(new_n966), .B2(new_n786), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(G1353gat));
  OR3_X1    g779(.A1(new_n962), .A2(G211gat), .A3(new_n608), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n964), .A2(new_n607), .A3(new_n903), .A4(new_n965), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n966), .B2(new_n633), .ZN(new_n987));
  OR3_X1    g786(.A1(new_n962), .A2(G218gat), .A3(new_n633), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1355gat));
endmodule


