//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(KEYINPUT69), .A3(G101), .A4(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(G137), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n461), .B2(new_n462), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n463), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G126), .A3(G2105), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n464), .A2(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(G543), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT70), .B1(new_n497), .B2(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n495), .A3(KEYINPUT6), .ZN(new_n500));
  AOI211_X1 g075(.A(new_n494), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G50), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(new_n494), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT71), .B(G88), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n502), .A2(new_n509), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  AND2_X1   g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n501), .A2(G51), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n498), .A2(new_n500), .ZN(new_n521));
  INV_X1    g096(.A(new_n496), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n521), .A2(G89), .A3(new_n522), .A4(new_n514), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT72), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  XOR2_X1   g104(.A(KEYINPUT73), .B(G52), .Z(new_n530));
  NAND3_X1  g105(.A1(new_n510), .A2(G543), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n510), .A2(G90), .A3(new_n514), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n512), .B2(new_n513), .ZN(new_n534));
  AND2_X1   g109(.A1(G77), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND4_X1  g113(.A1(new_n521), .A2(G43), .A3(G543), .A4(new_n522), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n521), .A2(G81), .A3(new_n522), .A4(new_n514), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI211_X1 g118(.A(KEYINPUT74), .B(new_n542), .C1(new_n506), .C2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n506), .B2(new_n543), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n495), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n541), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n512), .B2(new_n513), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(KEYINPUT75), .A2(G78), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n521), .A2(G91), .A3(new_n522), .A4(new_n514), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AND2_X1   g138(.A1(G53), .A2(G543), .ZN(new_n564));
  AND4_X1   g139(.A1(new_n563), .A2(new_n521), .A3(new_n522), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n510), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n561), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(G299));
  NAND3_X1  g142(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n510), .A2(G87), .A3(new_n514), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n501), .A2(G48), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n510), .A2(G86), .A3(new_n514), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n506), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(G305));
  NAND3_X1  g153(.A1(new_n510), .A2(G85), .A3(new_n514), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n510), .A2(G47), .A3(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n495), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT76), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n581), .A2(new_n495), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n584), .A2(new_n585), .A3(new_n579), .A4(new_n580), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n521), .A2(G92), .A3(new_n522), .A4(new_n514), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G66), .B1(new_n504), .B2(new_n505), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n495), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n501), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  OR3_X1    g177(.A1(G168), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT77), .B1(G168), .B2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n561), .A2(new_n562), .ZN(new_n605));
  INV_X1    g180(.A(new_n566), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n510), .A2(new_n563), .A3(new_n564), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n603), .B(new_n604), .C1(G868), .C2(new_n608), .ZN(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n599), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n545), .A2(new_n546), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n613), .A2(G651), .A3(new_n544), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n614), .A2(new_n539), .A3(new_n540), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n602), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n598), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g194(.A(G2104), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G2105), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n483), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n463), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n464), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n477), .A2(KEYINPUT79), .A3(G123), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT79), .B1(new_n477), .B2(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(G2096), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n626), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n638), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n649), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT17), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n657), .B1(new_n656), .B2(new_n654), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n655), .B2(new_n656), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n656), .A2(new_n654), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(new_n657), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(KEYINPUT84), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g258(.A(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT85), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT86), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n690), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n681), .B(new_n682), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n687), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n691), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n672), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n697), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n696), .A2(new_n687), .A3(new_n695), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n693), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n671), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(G171), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G5), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G1961), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G32), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n621), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n477), .A2(G129), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT27), .B(G1996), .Z(new_n721));
  AOI22_X1  g296(.A1(new_n710), .A2(new_n711), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G34), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT24), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(KEYINPUT24), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(KEYINPUT94), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT94), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n474), .B2(new_n712), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT95), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n722), .B1(new_n729), .B2(G2084), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT98), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n712), .A2(G33), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n463), .A2(G139), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n483), .A2(G127), .ZN(new_n738));
  INV_X1    g313(.A(G115), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n620), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n737), .B1(G2105), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n732), .B1(new_n741), .B2(new_n712), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G2072), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT93), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n712), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n712), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT96), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT30), .B2(new_n751), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n753), .C1(new_n632), .C2(new_n712), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n742), .B2(G2072), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n744), .A2(new_n748), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n463), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n477), .A2(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n464), .A2(G116), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n712), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n708), .A2(G20), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n608), .B2(new_n708), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1956), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n756), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n708), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n599), .B2(new_n708), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT90), .B(G1348), .Z(new_n776));
  XOR2_X1   g351(.A(new_n775), .B(new_n776), .Z(new_n777));
  NOR2_X1   g352(.A1(new_n710), .A2(new_n711), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n729), .A2(G2084), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT29), .B(G2090), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n720), .B2(new_n721), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G19), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n548), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1341), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n708), .A2(G21), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G286), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1966), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT97), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n789), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n731), .A2(new_n773), .A3(new_n785), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G6), .A2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1981), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n708), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n708), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT88), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT88), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n708), .A2(G22), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT89), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n708), .ZN(new_n813));
  INV_X1    g388(.A(G1971), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n803), .A2(new_n816), .A3(KEYINPUT34), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT34), .B1(new_n803), .B2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(G290), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G16), .B2(G24), .ZN(new_n821));
  INV_X1    g396(.A(G1986), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(G25), .A2(G29), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n463), .A2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n477), .A2(G119), .ZN(new_n827));
  OR2_X1    g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT87), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n823), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n817), .A2(new_n818), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n798), .B1(new_n838), .B2(new_n839), .ZN(G311));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  INV_X1    g416(.A(new_n798), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(G150));
  NAND4_X1  g418(.A1(new_n521), .A2(G55), .A3(G543), .A4(new_n522), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n521), .A2(G93), .A3(new_n522), .A4(new_n514), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n512), .B2(new_n513), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(KEYINPUT100), .B(new_n850), .C1(new_n506), .C2(new_n848), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(G651), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n846), .A2(KEYINPUT101), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n615), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n548), .A2(KEYINPUT101), .A3(new_n854), .A4(new_n846), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n599), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n855), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(G162), .B(new_n474), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n632), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n490), .A2(new_n492), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n484), .A2(new_n486), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n761), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n477), .A2(G130), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  INV_X1    g455(.A(G118), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(G2105), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n463), .A2(G142), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n879), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n877), .A2(new_n885), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n741), .B(new_n718), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n623), .B(new_n830), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n741), .B(new_n719), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n890), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n887), .A2(new_n888), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n887), .A2(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n873), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(new_n888), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n895), .A3(new_n872), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g480(.A1(new_n598), .A2(new_n608), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n565), .A2(new_n566), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n593), .B(new_n597), .C1(new_n907), .C2(new_n605), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(KEYINPUT104), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n599), .A2(new_n910), .A3(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n617), .A2(KEYINPUT103), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n617), .A2(KEYINPUT103), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(new_n861), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n915), .B1(new_n860), .B2(new_n859), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n906), .A2(new_n921), .A3(new_n908), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(new_n861), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n846), .A2(KEYINPUT101), .A3(new_n854), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT101), .B1(new_n846), .B2(new_n854), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(new_n548), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n615), .A2(new_n855), .A3(new_n856), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n914), .A3(new_n915), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n919), .A2(new_n931), .A3(KEYINPUT105), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n923), .A2(new_n924), .A3(new_n933), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g512(.A1(G303), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT106), .A4(new_n516), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n819), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(G290), .A2(new_n938), .A3(new_n939), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G305), .B(G288), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n932), .A2(new_n934), .A3(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n936), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n936), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n855), .A2(new_n602), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(G295));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n955), .ZN(G331));
  NAND2_X1  g532(.A1(G286), .A2(G301), .ZN(new_n958));
  OAI211_X1 g533(.A(G171), .B(new_n520), .C1(new_n526), .C2(new_n527), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n927), .B2(new_n928), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n859), .A2(new_n860), .A3(new_n958), .A4(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n929), .A2(KEYINPUT108), .A3(new_n958), .A4(new_n959), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n912), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n912), .A2(new_n921), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n906), .A2(new_n908), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT41), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n949), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n923), .A2(new_n964), .A3(new_n965), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n913), .A2(new_n963), .A3(new_n961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n948), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n899), .A4(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(new_n948), .A3(new_n975), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n948), .B1(new_n974), .B2(new_n975), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(new_n979), .A3(G37), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(new_n899), .A3(new_n976), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n973), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(KEYINPUT109), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n876), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n874), .B2(new_n875), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n469), .A2(new_n473), .A3(G40), .ZN(new_n998));
  OR3_X1    g573(.A1(new_n993), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n819), .A2(new_n822), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n718), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2067), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n761), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n831), .A2(new_n833), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n831), .A2(new_n833), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1003), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  INV_X1    g590(.A(new_n998), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1015), .B(new_n1016), .C1(new_n995), .C2(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1020), .B2(new_n1016), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n793), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G2084), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n876), .A2(new_n1025), .A3(new_n991), .ZN(new_n1026));
  AND4_X1   g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1016), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(G168), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1016), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT117), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1018), .A3(new_n1017), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1027), .B1(new_n1036), .B2(new_n793), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1033), .B1(new_n1037), .B2(G168), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT112), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n998), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n994), .C1(G164), .C2(G1384), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n747), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n998), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1026), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1043), .A2(new_n1048), .B1(new_n1050), .B2(new_n711), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1043), .A2(G2078), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1045), .B(new_n1052), .C1(new_n993), .C2(new_n997), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1051), .A2(G301), .A3(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1035), .A2(new_n1018), .A3(new_n1017), .A4(new_n1052), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1042), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G303), .A2(G8), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1058), .B(KEYINPUT55), .Z(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1024), .A2(new_n1016), .A3(new_n1026), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n814), .A2(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1058), .B(KEYINPUT55), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1016), .B1(new_n995), .B2(new_n1025), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1026), .A2(KEYINPUT116), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n995), .A2(new_n1069), .A3(new_n1025), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(new_n1063), .B1(new_n1061), .B2(new_n814), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1072), .B2(new_n1033), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1033), .B1(new_n995), .B2(new_n1016), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n568), .A2(new_n569), .A3(G1976), .A4(new_n570), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT114), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1080), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n995), .A2(new_n1016), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G8), .A3(new_n1075), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(KEYINPUT113), .A3(new_n1075), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(KEYINPUT52), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  INV_X1    g664(.A(G1981), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n577), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G305), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G305), .A2(new_n1092), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1095), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1098), .A3(new_n1074), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1082), .A2(new_n1088), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1065), .A2(new_n1073), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1051), .A2(G301), .A3(new_n1055), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1102), .B(KEYINPUT54), .C1(new_n1103), .C2(G301), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1041), .A2(new_n1057), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1070), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1069), .B1(new_n995), .B2(new_n1025), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1049), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT118), .B(G1956), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1050), .A2(new_n776), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n995), .A2(new_n1016), .A3(new_n1007), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n598), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1116), .B1(new_n1071), .B2(new_n1109), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1113), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1117), .A2(new_n1125), .A3(KEYINPUT61), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1117), .A2(new_n1125), .A3(KEYINPUT123), .A4(KEYINPUT61), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1044), .A2(new_n1045), .A3(new_n1005), .A4(new_n1047), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  AOI22_X1  g709(.A1(new_n1131), .A2(new_n1132), .B1(new_n1083), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n615), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1119), .A2(new_n1121), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT61), .B1(new_n1118), .B2(KEYINPUT122), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1117), .A2(new_n1125), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1130), .A2(new_n1138), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1105), .B1(new_n1123), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1031), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1039), .B1(new_n1038), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1030), .A2(KEYINPUT51), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT62), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1032), .A2(new_n1155), .A3(new_n1040), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1056), .A2(new_n1065), .A3(new_n1073), .A4(new_n1100), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1074), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1099), .A2(new_n1076), .A3(new_n805), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n800), .A2(new_n1090), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(G286), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1033), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1100), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1165), .B2(KEYINPUT63), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(G8), .A4(G168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1061), .A2(new_n814), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1049), .B(new_n1063), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1059), .B1(new_n1172), .B2(G8), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1065), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1100), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1166), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1158), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1014), .B1(new_n1150), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1008), .B(new_n719), .C1(new_n1179), .C2(G1996), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1003), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1000), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1179), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1182), .B2(new_n1179), .ZN(new_n1185));
  OAI211_X1 g760(.A(KEYINPUT47), .B(new_n1181), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1181), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT47), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1190), .A2(new_n1009), .B1(G2067), .B2(new_n761), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1003), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT124), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(KEYINPUT126), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT48), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1012), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1002), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1003), .A2(KEYINPUT48), .A3(new_n1012), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1003), .A2(new_n1200), .A3(new_n1011), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  AND4_X1   g777(.A1(new_n1186), .A2(new_n1189), .A3(new_n1193), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1178), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g779(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n1206), .A2(new_n706), .A3(new_n904), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n974), .A2(new_n975), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(new_n949), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n1209), .A2(new_n899), .A3(new_n976), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1210), .A2(KEYINPUT43), .ZN(new_n1211));
  AOI211_X1 g785(.A(KEYINPUT127), .B(new_n1207), .C1(new_n1211), .C2(new_n977), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1207), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n981), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1212), .A2(new_n1215), .ZN(G308));
  INV_X1    g790(.A(new_n977), .ZN(new_n1217));
  AOI21_X1  g791(.A(G37), .B1(new_n1208), .B2(new_n949), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n973), .B1(new_n1218), .B2(new_n976), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1214), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n1220), .A2(KEYINPUT127), .ZN(new_n1221));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1222), .ZN(G225));
endmodule


