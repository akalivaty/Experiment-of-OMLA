//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT29), .ZN(new_n210));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT76), .B(G155gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n212), .B1(new_n222), .B2(G162gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n211), .A2(new_n216), .A3(new_n218), .A4(new_n213), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n220), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(G22gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(G78gat), .B(G106gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT31), .B(G50gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G22gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n231), .B1(KEYINPUT80), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(G22gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n237), .B(KEYINPUT79), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT71), .ZN(new_n247));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n257), .A3(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT26), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n266), .B(KEYINPUT65), .C1(new_n248), .C2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  INV_X1    g069(.A(new_n248), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n272), .A3(new_n254), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  INV_X1    g074(.A(G190gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G183gat), .ZN(new_n281));
  AND4_X1   g080(.A1(new_n274), .A2(new_n279), .A3(new_n281), .A4(new_n276), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n273), .B1(new_n283), .B2(KEYINPUT28), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n277), .B2(new_n282), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT66), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n268), .A2(new_n272), .A3(new_n254), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n279), .A2(new_n281), .A3(new_n276), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT64), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT28), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT66), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n262), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n247), .B1(new_n295), .B2(new_n210), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n286), .A2(new_n288), .A3(new_n292), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n246), .B1(new_n297), .B2(new_n262), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n208), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n298), .B(KEYINPUT72), .ZN(new_n304));
  INV_X1    g103(.A(new_n247), .ZN(new_n305));
  INV_X1    g104(.A(new_n262), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n308), .B2(new_n293), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n305), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n209), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n262), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n210), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n295), .A2(new_n247), .B1(new_n246), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n209), .ZN(new_n316));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n312), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n301), .A2(new_n302), .B1(new_n209), .B2(new_n315), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n312), .A4(new_n319), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n316), .B1(new_n311), .B2(KEYINPUT73), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n302), .B(new_n209), .C1(new_n304), .C2(new_n310), .ZN(new_n328));
  INV_X1    g127(.A(new_n319), .ZN(new_n329));
  NOR4_X1   g128(.A1(new_n327), .A2(new_n328), .A3(new_n322), .A4(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n319), .B1(new_n323), .B2(new_n312), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  XOR2_X1   g133(.A(G127gat), .B(G134gat), .Z(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(KEYINPUT1), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT67), .B(G113gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(G120gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n348));
  OAI21_X1  g147(.A(G162gat), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n350));
  AND4_X1   g149(.A1(new_n216), .A2(new_n211), .A3(new_n218), .A4(new_n213), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n350), .A2(new_n351), .B1(new_n219), .B2(new_n214), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n346), .B1(new_n352), .B2(new_n221), .ZN(new_n353));
  INV_X1    g152(.A(new_n225), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n334), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n225), .A4(new_n346), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n341), .A2(G120gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n339), .ZN(new_n362));
  INV_X1    g161(.A(new_n345), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n338), .A2(G113gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n344), .B1(new_n340), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n362), .A2(new_n363), .B1(new_n365), .B2(new_n335), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n346), .B2(new_n227), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n355), .B2(new_n357), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n359), .A4(new_n360), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n366), .A2(new_n352), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n346), .A2(new_n227), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT5), .B1(new_n380), .B2(new_n360), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n374), .B2(new_n360), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n382), .B1(new_n373), .B2(new_n376), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT82), .B1(new_n392), .B2(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  OR3_X1    g194(.A1(new_n374), .A2(new_n395), .A3(new_n360), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n374), .B2(new_n360), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT39), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n380), .B2(new_n360), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n389), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT40), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT40), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n400), .A2(new_n405), .A3(new_n389), .A4(new_n402), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n245), .B1(new_n333), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n389), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT6), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n392), .B2(new_n389), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n411), .A3(new_n393), .ZN(new_n412));
  AND4_X1   g211(.A1(new_n410), .A2(new_n412), .A3(new_n321), .A4(new_n325), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n303), .A2(new_n312), .A3(new_n414), .A4(new_n316), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n323), .A2(KEYINPUT84), .A3(new_n414), .A4(new_n312), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n319), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n315), .B2(new_n208), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n296), .A2(new_n300), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n208), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n420), .B(KEYINPUT83), .C1(new_n208), .C2(new_n421), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n413), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n323), .A2(new_n312), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n408), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n308), .A2(new_n293), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n366), .B1(new_n442), .B2(new_n262), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n346), .B(new_n306), .C1(new_n308), .C2(new_n293), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n366), .B(new_n262), .C1(new_n287), .C2(new_n294), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT68), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT32), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n440), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n295), .A2(new_n346), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n309), .A2(new_n445), .A3(new_n366), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(new_n453), .A3(new_n441), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT32), .B1(new_n439), .B2(new_n450), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n448), .A2(new_n453), .A3(new_n454), .ZN(new_n459));
  INV_X1    g258(.A(new_n441), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n452), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n446), .A2(new_n456), .A3(new_n441), .A4(new_n448), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  INV_X1    g266(.A(new_n451), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n439), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT69), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT69), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n461), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n457), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n436), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n463), .A2(KEYINPUT36), .A3(new_n470), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT74), .B1(new_n330), .B2(new_n331), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n326), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n323), .A2(KEYINPUT30), .A3(new_n312), .A4(new_n319), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n327), .A2(new_n328), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n319), .ZN(new_n485));
  INV_X1    g284(.A(new_n411), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n410), .B1(new_n486), .B2(new_n409), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n245), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT70), .B(new_n436), .C1(new_n471), .C2(new_n474), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n479), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI221_X4 g290(.A(new_n319), .B1(new_n430), .B2(KEYINPUT37), .C1(new_n417), .C2(new_n418), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n413), .B(new_n427), .C1(new_n492), .C2(new_n429), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT85), .A3(new_n408), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n435), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n481), .A2(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n463), .A2(new_n470), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n245), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n471), .A2(new_n474), .ZN(new_n501));
  INV_X1    g300(.A(new_n333), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n245), .A2(KEYINPUT35), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n412), .A2(new_n410), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n495), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(KEYINPUT41), .ZN(new_n509));
  XNOR2_X1  g308(.A(G134gat), .B(G162gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT98), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT99), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT15), .B1(new_n515), .B2(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G50gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(G43gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT87), .B(G29gat), .Z(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT88), .A3(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT87), .B(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT89), .B1(new_n517), .B2(G43gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G43gat), .B2(new_n517), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT15), .B1(new_n518), .B2(KEYINPUT89), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n519), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n519), .B2(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT92), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n538));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G99gat), .B(G106gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n537), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n548), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(KEYINPUT41), .B2(new_n508), .ZN(new_n552));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n511), .A2(KEYINPUT98), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n550), .B2(new_n552), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n514), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(new_n555), .A3(new_n554), .A4(new_n513), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n217), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(G57gat), .ZN(new_n569));
  INV_X1    g368(.A(G57gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(KEYINPUT93), .A3(G64gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n571), .C1(new_n570), .C2(G64gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n574), .B(new_n581), .C1(new_n576), .C2(new_n580), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n575), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT96), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G231gat), .ZN(new_n592));
  INV_X1    g391(.A(G233gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G127gat), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n589), .B(new_n590), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(KEYINPUT90), .A2(G1gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(KEYINPUT90), .A2(G1gat), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT16), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT91), .ZN(new_n603));
  XNOR2_X1  g402(.A(G15gat), .B(G22gat), .ZN(new_n604));
  MUX2_X1   g403(.A(G1gat), .B(new_n603), .S(new_n604), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G8gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n588), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(KEYINPUT21), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n599), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G127gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n614), .B2(new_n598), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n566), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n599), .B2(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n612), .A3(new_n598), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n565), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n561), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n547), .B1(new_n586), .B2(new_n588), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n548), .B1(new_n582), .B2(new_n584), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT100), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT101), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n621), .B2(new_n622), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n626), .ZN(new_n638));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n606), .A2(new_n535), .ZN(new_n643));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n606), .A2(new_n538), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(new_n644), .C1(new_n537), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n606), .B(new_n535), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n644), .B(KEYINPUT13), .Z(new_n649));
  AOI22_X1  g448(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n537), .A2(new_n645), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n644), .A4(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G169gat), .B(G197gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n650), .A2(new_n652), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n507), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n487), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g468(.A1(new_n666), .A2(new_n333), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n674));
  INV_X1    g473(.A(G8gat), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n670), .ZN(G1325gat));
  AOI21_X1  g475(.A(G15gat), .B1(new_n666), .B2(new_n501), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n479), .A2(new_n490), .ZN(new_n679));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT103), .Z(new_n682));
  AOI21_X1  g481(.A(new_n678), .B1(new_n666), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n245), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  AND3_X1   g485(.A1(new_n493), .A2(KEYINPUT85), .A3(new_n408), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT85), .B1(new_n493), .B2(new_n408), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n479), .A2(new_n489), .A3(new_n490), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n506), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n561), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n616), .A2(new_n619), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n637), .A2(new_n640), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n694), .A2(new_n664), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n520), .B1(new_n697), .B2(new_n487), .ZN(new_n698));
  INV_X1    g497(.A(new_n561), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n495), .B2(new_n506), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n667), .A3(new_n523), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(G1328gat));
  OAI21_X1  g503(.A(G36gat), .B1(new_n697), .B2(new_n502), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(new_n524), .A3(new_n333), .ZN(new_n706));
  AND2_X1   g505(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n705), .B(new_n709), .C1(new_n707), .C2(new_n706), .ZN(G1329gat));
  OR2_X1    g509(.A1(new_n679), .A2(new_n515), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n701), .A2(new_n501), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n697), .A2(new_n711), .B1(G43gat), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g513(.A(new_n245), .ZN(new_n715));
  OAI21_X1  g514(.A(G50gat), .B1(new_n697), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n245), .A2(new_n517), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT105), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  NAND4_X1  g523(.A1(new_n507), .A2(new_n664), .A3(new_n620), .A4(new_n695), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n487), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n570), .ZN(G1332gat));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n502), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  AND2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n728), .B2(new_n729), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n725), .B2(new_n679), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n501), .A2(new_n578), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n725), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g535(.A1(new_n725), .A2(new_n715), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT106), .B(G78gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1335gat));
  NAND3_X1  g538(.A1(new_n695), .A2(new_n667), .A3(new_n542), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n694), .A2(new_n663), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n692), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n700), .A2(KEYINPUT107), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n700), .B2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n744), .B(new_n699), .C1(new_n495), .C2(new_n506), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n741), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n692), .A2(new_n744), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n742), .A4(new_n746), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT108), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n740), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n743), .A2(new_n641), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n693), .A2(new_n667), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G85gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT109), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n740), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT108), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT108), .B1(new_n753), .B2(new_n755), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n760), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n693), .A2(new_n333), .A3(new_n758), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n747), .A2(new_n751), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n333), .A2(new_n695), .A3(new_n543), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n771), .B(new_n776), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1337gat));
  INV_X1    g577(.A(new_n501), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n779), .A2(G99gat), .A3(new_n641), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n764), .B2(new_n765), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n693), .A2(new_n758), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n782), .B2(new_n679), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1338gat));
  NAND3_X1  g583(.A1(new_n693), .A2(new_n245), .A3(new_n758), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n641), .A2(new_n715), .A3(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n772), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n786), .B(new_n790), .C1(new_n772), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1339gat));
  NAND3_X1  g591(.A1(new_n629), .A2(new_n625), .A3(new_n630), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n636), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n663), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n637), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n644), .B1(new_n651), .B2(new_n643), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n648), .A2(new_n649), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n658), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n662), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n801), .A2(new_n803), .B1(new_n641), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n699), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n637), .A2(new_n802), .ZN(new_n810));
  INV_X1    g609(.A(new_n807), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n810), .A2(new_n561), .A3(new_n811), .A4(new_n800), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n694), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n620), .A2(new_n664), .A3(new_n641), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n245), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n333), .A2(new_n487), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n501), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n664), .ZN(new_n822));
  INV_X1    g621(.A(new_n812), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n699), .B2(new_n808), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n814), .B1(new_n824), .B2(new_n694), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n667), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n245), .A3(new_n497), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n502), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n663), .A2(new_n341), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  OAI21_X1  g629(.A(new_n338), .B1(new_n828), .B2(new_n641), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n820), .A2(G120gat), .A3(new_n695), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT110), .Z(G1341gat));
  INV_X1    g633(.A(new_n694), .ZN(new_n835));
  OAI21_X1  g634(.A(G127gat), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n694), .A2(new_n596), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n828), .B2(new_n837), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n699), .A2(G134gat), .A3(new_n333), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n827), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT111), .Z(new_n842));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n561), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n843), .B2(G134gat), .ZN(new_n844));
  INV_X1    g643(.A(new_n840), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n667), .A2(new_n825), .A3(new_n245), .A4(new_n679), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n502), .ZN(new_n851));
  INV_X1    g650(.A(G141gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n663), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n679), .A2(new_n818), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n660), .A2(new_n662), .B1(new_n798), .B2(new_n799), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n856), .A2(new_n810), .B1(new_n695), .B2(new_n811), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n561), .B1(new_n857), .B2(KEYINPUT113), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n808), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n823), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n814), .B1(new_n861), .B2(new_n694), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n245), .ZN(new_n863));
  XOR2_X1   g662(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n816), .B2(new_n715), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n855), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n852), .B1(new_n866), .B2(new_n663), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n853), .A2(new_n333), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n848), .B2(new_n868), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n854), .A2(new_n867), .B1(new_n869), .B2(new_n847), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n641), .A2(G148gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n502), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  INV_X1    g672(.A(new_n855), .ZN(new_n874));
  INV_X1    g673(.A(new_n864), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n245), .B(new_n875), .C1(new_n813), .C2(new_n815), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT115), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n825), .A2(new_n878), .A3(new_n245), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n814), .B(KEYINPUT116), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n861), .B2(new_n694), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n245), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n695), .B(new_n874), .C1(new_n880), .C2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n873), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n873), .A2(G148gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n866), .B2(new_n695), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n872), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n872), .B(new_n890), .C1(new_n885), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1345gat));
  INV_X1    g691(.A(new_n866), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n222), .B1(new_n893), .B2(new_n835), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n835), .A2(new_n222), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n851), .B2(new_n895), .ZN(G1346gat));
  NAND4_X1  g695(.A1(new_n850), .A2(new_n215), .A3(new_n502), .A4(new_n561), .ZN(new_n897));
  OAI21_X1  g696(.A(G162gat), .B1(new_n893), .B2(new_n699), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NAND3_X1  g698(.A1(new_n501), .A2(new_n487), .A3(new_n333), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT120), .Z(new_n901));
  NAND3_X1  g700(.A1(new_n825), .A2(new_n901), .A3(new_n715), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n264), .A3(new_n664), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n816), .A2(new_n667), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n498), .A2(new_n333), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT118), .Z(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n663), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(new_n264), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n265), .A3(new_n695), .ZN(new_n911));
  OAI21_X1  g710(.A(G176gat), .B1(new_n902), .B2(new_n641), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  NAND4_X1  g712(.A1(new_n817), .A2(KEYINPUT122), .A3(new_n694), .A4(new_n901), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n902), .B2(new_n835), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n916), .A3(G183gat), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n694), .A2(new_n275), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n825), .A2(new_n487), .A3(new_n906), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  AND2_X1   g721(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n917), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n922), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n908), .A2(new_n276), .A3(new_n561), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n902), .B2(new_n699), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n679), .A2(new_n245), .A3(new_n333), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n904), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n663), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n880), .A2(new_n883), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n679), .A2(new_n487), .A3(new_n333), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT127), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n663), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n946), .B2(new_n938), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n941), .A2(new_n695), .A3(new_n943), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G204gat), .ZN(new_n949));
  INV_X1    g748(.A(G204gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n950), .A3(new_n695), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n203), .A3(new_n694), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n694), .A3(new_n943), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n937), .A2(new_n204), .A3(new_n561), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n561), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n962), .B2(new_n204), .ZN(G1355gat));
endmodule


