//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n191), .B2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G119), .ZN(new_n193));
  MUX2_X1   g007(.A(KEYINPUT23), .B(new_n192), .S(new_n193), .Z(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  OAI22_X1  g010(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n201), .B(new_n203), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n194), .A2(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n196), .A2(new_n195), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(KEYINPUT76), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(KEYINPUT76), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n190), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n190), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n210), .B2(KEYINPUT76), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OR3_X1    g030(.A1(new_n216), .A2(KEYINPUT25), .A3(G902), .ZN(new_n217));
  INV_X1    g031(.A(G217), .ZN(new_n218));
  INV_X1    g032(.A(G902), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(G234), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT25), .B1(new_n216), .B2(G902), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n220), .A2(G902), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT77), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n227), .B(KEYINPUT11), .C1(new_n228), .C2(G137), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  OAI211_X1 g045(.A(G134), .B(new_n230), .C1(new_n231), .C2(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n230), .A2(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n236), .A2(new_n237), .B1(KEYINPUT64), .B2(new_n231), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n233), .A2(new_n238), .A3(new_n241), .A4(new_n235), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(KEYINPUT66), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n244), .A3(G131), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT0), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n191), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT0), .B(G128), .Z(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n243), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n228), .A2(G137), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n242), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n191), .A2(new_n203), .A3(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n246), .B2(new_n256), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n203), .A2(G143), .ZN(new_n262));
  AND4_X1   g076(.A1(KEYINPUT67), .A2(new_n256), .A3(new_n262), .A4(new_n258), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n255), .B(new_n260), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n256), .A2(new_n262), .A3(new_n258), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n246), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n259), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n274), .B1(new_n279), .B2(new_n255), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n254), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n251), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n281), .A2(new_n284), .A3(KEYINPUT30), .A4(new_n251), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G119), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n289));
  INV_X1    g103(.A(G119), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(G116), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(KEYINPUT69), .A3(G119), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT2), .B(G113), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n293), .B2(new_n294), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n272), .A2(new_n286), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n295), .B(KEYINPUT70), .ZN(new_n300));
  INV_X1    g114(.A(new_n293), .ZN(new_n301));
  INV_X1    g115(.A(new_n294), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n281), .A3(new_n251), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n188), .A3(G210), .ZN(new_n306));
  INV_X1    g120(.A(G101), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n308), .B(new_n309), .Z(new_n310));
  NAND3_X1  g124(.A1(new_n299), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT31), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT31), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n299), .A2(new_n313), .A3(new_n304), .A4(new_n310), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n266), .A2(new_n298), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n304), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT73), .B1(new_n281), .B2(new_n251), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n281), .A2(KEYINPUT73), .A3(new_n251), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n303), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n315), .B1(new_n323), .B2(new_n310), .ZN(new_n324));
  INV_X1    g138(.A(new_n310), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n303), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n316), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT74), .B(new_n325), .C1(new_n328), .C2(new_n318), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n312), .A2(new_n314), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G472), .A2(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT32), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(new_n304), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n269), .A2(new_n271), .B1(new_n283), .B2(new_n285), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n298), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n325), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n310), .B1(new_n328), .B2(new_n318), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n303), .B1(new_n251), .B2(new_n281), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT28), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n219), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G472), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n334), .A2(new_n335), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n334), .A2(KEYINPUT75), .A3(new_n335), .A4(new_n347), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n226), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G221), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT9), .B(G234), .Z(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n219), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G469), .ZN(new_n357));
  XNOR2_X1  g171(.A(G110), .B(G140), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n188), .A2(G227), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g174(.A(KEYINPUT12), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n362), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G107), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n366), .A3(new_n307), .A4(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(G104), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n307), .B1(new_n372), .B2(new_n367), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n264), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n373), .B1(new_n369), .B2(new_n370), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n264), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n377), .A2(new_n380), .B1(new_n376), .B2(new_n375), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n243), .A2(new_n245), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n361), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n380), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n379), .B1(new_n378), .B2(new_n264), .ZN(new_n385));
  OAI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(new_n264), .B2(new_n378), .ZN(new_n386));
  INV_X1    g200(.A(new_n382), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT12), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n384), .B2(new_n385), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n371), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n393), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n250), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n378), .B(KEYINPUT10), .C1(new_n273), .C2(new_n280), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n391), .A2(new_n399), .A3(new_n382), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n360), .B1(new_n389), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n391), .A2(new_n399), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n387), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n401), .A3(new_n360), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(KEYINPUT81), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n402), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n357), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n360), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n388), .B2(new_n383), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n360), .B1(new_n405), .B2(new_n401), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n357), .B(new_n219), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n357), .A2(new_n219), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n396), .A2(new_n298), .A3(new_n397), .A4(new_n398), .ZN(new_n420));
  INV_X1    g234(.A(G113), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n288), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n301), .A2(new_n422), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n300), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n378), .ZN(new_n426));
  XOR2_X1   g240(.A(G110), .B(G122), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n264), .A2(new_n198), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n250), .A2(G125), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n188), .A2(G224), .B1(KEYINPUT83), .B2(KEYINPUT7), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(KEYINPUT83), .B2(KEYINPUT7), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n431), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n188), .A2(G224), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(KEYINPUT7), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n375), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n423), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n378), .B1(new_n300), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n427), .B(KEYINPUT8), .Z(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n429), .A2(new_n439), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n219), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n420), .A2(new_n426), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n427), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n436), .B(new_n437), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n455), .A3(new_n427), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n219), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n450), .A2(new_n457), .A3(new_n460), .A4(new_n458), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n305), .A2(new_n188), .A3(G214), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(G143), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n241), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT17), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n241), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n206), .B(new_n471), .C1(new_n472), .C2(KEYINPUT17), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(KEYINPUT18), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT18), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n475), .B2(new_n241), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n200), .B(new_n203), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G113), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n362), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n481), .A2(KEYINPUT87), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n481), .ZN(new_n486));
  INV_X1    g300(.A(G475), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT19), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n490));
  MUX2_X1   g304(.A(new_n489), .B(new_n490), .S(new_n200), .Z(new_n491));
  OAI211_X1 g305(.A(new_n472), .B(new_n202), .C1(G146), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n481), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n478), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n486), .A2(new_n487), .A3(new_n219), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n485), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n188), .A2(G952), .ZN(new_n501));
  NAND2_X1  g315(.A1(G234), .A2(G237), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT90), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(G902), .A3(G953), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G128), .B(G143), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n228), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT88), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n287), .A2(KEYINPUT14), .A3(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(G116), .B(G122), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(G107), .B(new_n511), .C1(new_n513), .C2(KEYINPUT14), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(G107), .B2(new_n513), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n228), .B(new_n516), .C1(KEYINPUT13), .C2(new_n508), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n512), .B(new_n365), .ZN(new_n518));
  INV_X1    g332(.A(new_n508), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(G134), .B2(new_n519), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n510), .A2(new_n515), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n354), .A2(G217), .A3(new_n188), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n219), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n526), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n500), .A2(new_n507), .A3(new_n534), .ZN(new_n535));
  AND4_X1   g349(.A1(new_n356), .A2(new_n419), .A3(new_n467), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n352), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT91), .B(G101), .Z(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(G3));
  NAND2_X1  g353(.A1(new_n330), .A2(new_n219), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G472), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n332), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n356), .B1(new_n411), .B2(new_n418), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n542), .A2(new_n226), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n467), .A2(new_n507), .ZN(new_n546));
  INV_X1    g360(.A(new_n522), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT33), .B1(new_n547), .B2(KEYINPUT93), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n524), .B2(new_n525), .ZN(new_n549));
  INV_X1    g363(.A(new_n525), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n523), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n527), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n527), .B(new_n219), .C1(new_n524), .C2(new_n525), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n527), .A2(new_n219), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n500), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n546), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n545), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT94), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT34), .B(G104), .Z(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(G6));
  INV_X1    g379(.A(new_n546), .ZN(new_n566));
  INV_X1    g380(.A(new_n498), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT95), .B1(new_n567), .B2(new_n496), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n496), .A2(KEYINPUT95), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND4_X1   g384(.A1(new_n485), .A2(new_n566), .A3(new_n533), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n545), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G107), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G9));
  NOR2_X1   g388(.A1(new_n214), .A2(KEYINPUT36), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n210), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n223), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n222), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n536), .A2(new_n332), .A3(new_n541), .A4(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT37), .B(G110), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G12));
  OAI21_X1  g395(.A(new_n504), .B1(G900), .B2(new_n506), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n485), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n533), .B(new_n583), .C1(new_n568), .C2(new_n569), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n586), .A2(new_n543), .A3(new_n466), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n330), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT32), .B1(new_n330), .B2(new_n331), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT75), .B1(new_n590), .B2(new_n347), .ZN(new_n591));
  INV_X1    g405(.A(new_n351), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n587), .B(new_n578), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G128), .ZN(G30));
  XOR2_X1   g408(.A(new_n582), .B(KEYINPUT39), .Z(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n419), .A2(new_n356), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n465), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n464), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n462), .A2(new_n463), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n499), .A2(new_n533), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n338), .A2(new_n325), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n336), .A2(new_n342), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n219), .B1(new_n611), .B2(new_n310), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n334), .A2(new_n335), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n578), .B1(new_n597), .B2(new_n598), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n601), .A2(new_n609), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G143), .ZN(G45));
  NAND2_X1  g431(.A1(new_n559), .A2(new_n582), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n543), .A2(new_n466), .A3(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n578), .B(new_n619), .C1(new_n591), .C2(new_n592), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G146), .ZN(G48));
  OR2_X1    g435(.A1(new_n413), .A2(new_n414), .ZN(new_n622));
  NAND2_X1  g436(.A1(KEYINPUT99), .A2(G469), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n219), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n413), .A2(new_n414), .ZN(new_n625));
  OAI211_X1 g439(.A(KEYINPUT99), .B(G469), .C1(new_n625), .C2(G902), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n624), .A2(new_n626), .A3(new_n356), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n352), .A2(new_n561), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n352), .A2(new_n630), .A3(new_n561), .A4(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT41), .B(G113), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G15));
  AND2_X1   g448(.A1(new_n352), .A2(new_n627), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n571), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G116), .ZN(G18));
  NAND2_X1  g451(.A1(new_n350), .A2(new_n351), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n624), .A2(new_n626), .A3(new_n356), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n466), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n638), .A2(new_n535), .A3(new_n578), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT101), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n350), .A2(new_n351), .B1(new_n222), .B2(new_n577), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n535), .A4(new_n640), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(G119), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G21));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n541), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n327), .A2(new_n343), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n327), .B2(new_n343), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n655), .A3(new_n310), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n313), .B1(new_n338), .B2(new_n310), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n655), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n653), .A3(new_n325), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n312), .A3(KEYINPUT104), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n314), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n331), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n226), .A2(KEYINPUT106), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n222), .B2(new_n225), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n540), .A2(KEYINPUT105), .A3(G472), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n650), .A2(new_n663), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n669), .A2(new_n546), .A3(new_n608), .A4(new_n639), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(G122), .Z(G24));
  INV_X1    g485(.A(new_n331), .ZN(new_n672));
  INV_X1    g486(.A(new_n314), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n660), .A2(new_n312), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n651), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n675), .B2(new_n661), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT105), .B1(new_n540), .B2(G472), .ZN(new_n677));
  INV_X1    g491(.A(G472), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n649), .B(new_n678), .C1(new_n330), .C2(new_n219), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n618), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n578), .A3(new_n681), .A4(new_n640), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G125), .ZN(G27));
  NOR2_X1   g497(.A1(new_n409), .A2(new_n402), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n418), .B1(G469), .B2(new_n684), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n685), .A2(new_n464), .A3(new_n355), .A4(new_n600), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n618), .A2(KEYINPUT42), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n352), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n681), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n335), .A2(KEYINPUT107), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n330), .A2(new_n691), .A3(KEYINPUT32), .A4(new_n331), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n334), .A3(new_n347), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n667), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G131), .ZN(G33));
  INV_X1    g511(.A(new_n586), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n352), .A2(new_n698), .A3(new_n686), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G134), .ZN(G36));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n407), .A2(new_n701), .A3(new_n410), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n357), .B1(new_n684), .B2(KEYINPUT45), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n416), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n625), .A2(G469), .A3(G902), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n704), .B2(KEYINPUT46), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n355), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n596), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n558), .A2(KEYINPUT43), .A3(new_n499), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n500), .B2(new_n557), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n542), .A2(new_n578), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n709), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n464), .A2(new_n600), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n716), .B(new_n717), .C1(new_n710), .C2(new_n715), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G137), .ZN(G39));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT47), .B(new_n355), .C1(new_n705), .C2(new_n707), .ZN(new_n722));
  INV_X1    g536(.A(new_n717), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n618), .A4(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n350), .A3(new_n351), .A4(new_n226), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT108), .B(G140), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G42));
  NAND2_X1  g541(.A1(new_n624), .A2(new_n626), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT49), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n558), .A2(new_n499), .A3(new_n355), .A4(new_n600), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n667), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT109), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT110), .B1(new_n728), .B2(KEYINPUT49), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n728), .A2(KEYINPUT110), .A3(KEYINPUT49), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n614), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n607), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n578), .B1(new_n590), .B2(new_n613), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n466), .A2(new_n685), .A3(new_n608), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n356), .A3(new_n582), .A4(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n593), .A2(new_n620), .A3(new_n682), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT112), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n643), .B1(new_n587), .B2(new_n619), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n682), .A4(new_n739), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n741), .A2(KEYINPUT52), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(new_n741), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n670), .B1(new_n635), .B2(new_n571), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n560), .B1(new_n499), .B2(new_n534), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n544), .A2(new_n566), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n537), .A2(new_n579), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n632), .A2(new_n748), .A3(new_n646), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n650), .A2(new_n663), .A3(new_n578), .A4(new_n668), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n681), .A3(new_n686), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n717), .A2(new_n534), .A3(new_n583), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n419), .A2(new_n356), .A3(new_n570), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n638), .A2(new_n578), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n696), .A2(new_n699), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT53), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n688), .A2(new_n699), .A3(new_n759), .A4(new_n695), .ZN(new_n763));
  INV_X1    g577(.A(new_n755), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n629), .A2(new_n631), .B1(new_n642), .B2(new_n645), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n748), .A4(new_n751), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n740), .A2(KEYINPUT111), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n740), .B2(KEYINPUT111), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n767), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n762), .A2(new_n773), .A3(KEYINPUT54), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n747), .A2(KEYINPUT53), .A3(new_n761), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n772), .B1(new_n767), .B2(new_n771), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n504), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n714), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n669), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n627), .A2(new_n604), .A3(new_n600), .A4(new_n605), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT50), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n669), .A2(new_n782), .A3(new_n785), .A4(new_n780), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT114), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n780), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n680), .A2(new_n667), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n785), .B1(new_n789), .B2(new_n782), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(KEYINPUT50), .A3(new_n783), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n627), .A2(new_n717), .A3(new_n779), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n558), .A2(new_n500), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n794), .A2(new_n614), .A3(new_n226), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n714), .A2(new_n627), .A3(new_n717), .A4(new_n779), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n753), .A2(new_n797), .A3(KEYINPUT115), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n753), .B2(new_n797), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n787), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT116), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n356), .B1(new_n728), .B2(KEYINPUT113), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(KEYINPUT113), .B2(new_n728), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n721), .B2(new_n722), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n717), .A3(new_n781), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n787), .A2(new_n793), .A3(new_n807), .A4(new_n800), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n798), .A2(new_n799), .ZN(new_n812));
  INV_X1    g626(.A(new_n796), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n810), .B1(new_n790), .B2(new_n791), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n800), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n816), .A3(new_n806), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n812), .B2(new_n813), .ZN(new_n821));
  AOI211_X1 g635(.A(KEYINPUT117), .B(new_n796), .C1(new_n798), .C2(new_n799), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n816), .A4(new_n806), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n694), .A2(new_n827), .A3(new_n797), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n694), .B2(new_n797), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(KEYINPUT121), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(KEYINPUT48), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n781), .A2(new_n640), .ZN(new_n835));
  OR4_X1    g649(.A1(new_n226), .A2(new_n794), .A3(new_n614), .A4(new_n560), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT48), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n501), .B(KEYINPUT119), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n811), .A2(new_n826), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n774), .A2(new_n778), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(G952), .A2(G953), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n736), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT122), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n736), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(G75));
  NAND2_X1  g663(.A1(new_n747), .A2(new_n761), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n772), .ZN(new_n851));
  INV_X1    g665(.A(new_n773), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n219), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(G210), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n453), .A2(new_n456), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(new_n454), .ZN(new_n857));
  XOR2_X1   g671(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n854), .B2(new_n855), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n188), .A2(G952), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G51));
  NAND2_X1  g677(.A1(new_n417), .A2(KEYINPUT57), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n417), .A2(KEYINPUT57), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n775), .B1(new_n851), .B2(new_n852), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n774), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n622), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n853), .A2(new_n702), .A3(new_n703), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(G54));
  NAND3_X1  g684(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n486), .A2(new_n494), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n862), .ZN(G60));
  INV_X1    g689(.A(new_n862), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n556), .B(KEYINPUT59), .ZN(new_n877));
  INV_X1    g691(.A(new_n778), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n851), .A2(new_n852), .A3(new_n775), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n549), .A2(new_n552), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n866), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n877), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n881), .B2(new_n884), .ZN(G63));
  NAND2_X1  g699(.A1(G217), .A2(G902), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT60), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n851), .B2(new_n852), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n862), .B1(new_n888), .B2(new_n576), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n891));
  INV_X1    g705(.A(new_n887), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n762), .B2(new_n773), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n216), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n890), .A2(new_n891), .ZN(new_n897));
  INV_X1    g711(.A(new_n894), .ZN(new_n898));
  INV_X1    g712(.A(new_n576), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n876), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n895), .A2(new_n901), .ZN(G66));
  AOI21_X1  g716(.A(new_n188), .B1(new_n505), .B2(G224), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n752), .B2(new_n188), .ZN(new_n904));
  INV_X1    g718(.A(G898), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n856), .B1(new_n905), .B2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n904), .B(new_n906), .ZN(G69));
  NAND2_X1  g721(.A1(G900), .A2(G953), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n337), .B(new_n491), .Z(new_n909));
  AND2_X1   g723(.A1(new_n742), .A2(new_n682), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n696), .ZN(new_n911));
  INV_X1    g725(.A(new_n699), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n709), .A2(new_n694), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n466), .A2(new_n608), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n911), .A2(new_n725), .A3(new_n718), .A4(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n908), .B(new_n909), .C1(new_n916), .C2(G953), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n597), .A2(new_n723), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n352), .A2(new_n749), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n725), .A2(new_n718), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n910), .A2(new_n616), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT127), .Z(new_n927));
  AOI21_X1  g741(.A(G953), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n909), .B(KEYINPUT125), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G72));
  INV_X1    g746(.A(new_n339), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n933), .B(new_n610), .C1(new_n776), .C2(new_n777), .ZN(new_n934));
  NAND2_X1  g748(.A1(G472), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT63), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n916), .B2(new_n752), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n862), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n925), .A2(new_n927), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n936), .B1(new_n941), .B2(new_n752), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n610), .B2(new_n942), .ZN(G57));
endmodule


