//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(KEYINPUT83), .A3(G125), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n190), .A2(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n188), .A2(G143), .ZN(new_n202));
  OAI211_X1 g016(.A(G128), .B(new_n200), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n189), .B(new_n191), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(new_n199), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G224), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G953), .ZN(new_n211));
  XOR2_X1   g025(.A(new_n209), .B(new_n211), .Z(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G104), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(G107), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n215), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G104), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(new_n222), .B2(new_n220), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n225));
  AOI211_X1 g039(.A(new_n225), .B(new_n219), .C1(new_n222), .C2(new_n220), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT2), .B(G113), .Z(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n231), .B2(G116), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(G119), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n230), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n232), .B2(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n240), .B2(new_n237), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n239), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n247));
  XNOR2_X1  g061(.A(G104), .B(G107), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n225), .B1(new_n248), .B2(new_n219), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n229), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n215), .A2(new_n218), .A3(new_n220), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G101), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n242), .A2(new_n230), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n239), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(G101), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT79), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G122), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n242), .B(new_n230), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n255), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n252), .A2(new_n260), .A3(new_n261), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(KEYINPUT81), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n252), .A2(new_n260), .A3(new_n265), .ZN(new_n273));
  INV_X1    g087(.A(new_n261), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n274), .A3(new_n272), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n213), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n252), .A2(new_n265), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT82), .A3(new_n261), .A4(new_n260), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n266), .A2(new_n267), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT7), .B1(new_n210), .B2(G953), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n209), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n285), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n198), .A2(new_n199), .A3(new_n208), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(new_n245), .ZN(new_n291));
  OR3_X1    g105(.A1(new_n291), .A2(new_n227), .A3(new_n239), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n293));
  INV_X1    g107(.A(new_n227), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n246), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n243), .A2(new_n245), .ZN(new_n296));
  OAI211_X1 g110(.A(KEYINPUT85), .B(new_n227), .C1(new_n296), .C2(new_n239), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(new_n261), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n289), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n284), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n279), .A2(new_n280), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n280), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n273), .A2(new_n274), .A3(new_n272), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(new_n275), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n212), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n301), .B1(new_n268), .B2(new_n269), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n304), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(G953), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n315), .A2(G952), .ZN(new_n316));
  INV_X1    g130(.A(G234), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n310), .B(new_n315), .C1(G234), .C2(G237), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT21), .B(G898), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n314), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G221), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT9), .B(G234), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n310), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT74), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n227), .A2(new_n206), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n250), .A2(new_n205), .A3(new_n203), .A4(new_n221), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G134), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G137), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G137), .ZN(new_n337));
  INV_X1    g151(.A(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT11), .A3(G134), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n336), .A2(new_n339), .A3(new_n342), .A4(new_n337), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n333), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  INV_X1    g160(.A(new_n344), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n346), .B(new_n347), .C1(new_n331), .C2(new_n332), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT78), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n227), .A2(new_n206), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n250), .A2(new_n221), .B1(new_n205), .B2(new_n203), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n333), .A2(KEYINPUT12), .A3(new_n344), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n253), .A2(G101), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n195), .B1(new_n358), .B2(new_n254), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n332), .A2(new_n357), .B1(new_n359), .B2(new_n264), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n200), .A2(G128), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n193), .ZN(new_n363));
  INV_X1    g177(.A(new_n205), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n203), .A2(KEYINPUT65), .A3(new_n205), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n229), .A2(new_n367), .A3(KEYINPUT10), .A4(new_n251), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n344), .B(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G140), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n315), .A2(G227), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n349), .A2(new_n356), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n371), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n347), .B1(new_n360), .B2(new_n368), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G469), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n310), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n310), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n371), .A2(new_n375), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n371), .B1(new_n348), .B2(new_n345), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n384), .A2(new_n385), .B1(new_n386), .B2(new_n374), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n387), .B2(G469), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n330), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G128), .B(G143), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n335), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G116), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n234), .A2(G122), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n217), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n234), .A2(KEYINPUT14), .A3(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n394), .ZN(new_n397));
  OAI211_X1 g211(.A(G107), .B(new_n396), .C1(new_n397), .C2(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n217), .B1(new_n393), .B2(new_n394), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n395), .A3(KEYINPUT90), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n403));
  INV_X1    g217(.A(new_n395), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n400), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n190), .A2(G128), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n335), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n204), .A2(G143), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n413), .A3(new_n335), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n390), .A2(KEYINPUT92), .A3(new_n335), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n410), .A2(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n406), .A2(new_n418), .A3(KEYINPUT93), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT93), .B1(new_n406), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n399), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n327), .A2(new_n423), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n418), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n419), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n399), .A3(new_n424), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G478), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT94), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(G902), .B(new_n438), .C1(new_n426), .C2(new_n431), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G140), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G125), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n207), .A2(G140), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT16), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n207), .A2(G140), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n188), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n449), .A3(G146), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT71), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n454), .A3(new_n188), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AND4_X1   g270(.A1(G143), .A2(new_n318), .A3(new_n315), .A4(G214), .ZN(new_n457));
  NOR2_X1   g271(.A1(G237), .A2(G953), .ZN(new_n458));
  AOI21_X1  g272(.A(G143), .B1(new_n458), .B2(G214), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n318), .A2(new_n315), .A3(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n190), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(G143), .A3(G214), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n342), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n465), .A2(KEYINPUT17), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT17), .A3(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n457), .A2(new_n459), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n444), .A2(new_n445), .A3(new_n188), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n443), .A2(G125), .ZN(new_n473));
  OAI21_X1  g287(.A(G146), .B1(new_n447), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n470), .A2(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT86), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n478), .B(new_n471), .C1(new_n462), .C2(new_n463), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G113), .B(G122), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n214), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n453), .A2(new_n455), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n468), .B1(new_n465), .B2(KEYINPUT17), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n483), .B(new_n480), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G475), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT19), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT19), .B1(new_n444), .B2(new_n445), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n188), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n465), .A2(new_n452), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(KEYINPUT87), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n484), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT87), .B1(new_n480), .B2(new_n495), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT88), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n474), .A2(new_n472), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n462), .A2(new_n463), .A3(new_n471), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n478), .B1(new_n470), .B2(new_n471), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n467), .A2(KEYINPUT86), .A3(new_n476), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n465), .A2(new_n452), .A3(new_n494), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n484), .A3(new_n496), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n488), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n500), .A2(new_n501), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT20), .ZN(new_n515));
  NOR3_X1   g329(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT89), .B(new_n517), .C1(new_n511), .C2(new_n488), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n499), .B2(new_n516), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n491), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n389), .A2(new_n442), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n187), .B1(new_n325), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n442), .ZN(new_n525));
  INV_X1    g339(.A(new_n330), .ZN(new_n526));
  AOI211_X1 g340(.A(G469), .B(G902), .C1(new_n376), .C2(new_n379), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n385), .A2(new_n384), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n386), .A2(new_n374), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(G469), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n383), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n526), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n314), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n303), .B2(new_n312), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n534), .A2(KEYINPUT95), .A3(new_n536), .A4(new_n324), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n423), .B1(G234), .B2(new_n310), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT22), .B(G137), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n326), .A2(new_n317), .A3(G953), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n231), .A2(G128), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT69), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n231), .B2(G128), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT69), .B1(new_n231), .B2(G128), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT70), .B1(new_n549), .B2(G110), .ZN(new_n550));
  XNOR2_X1  g364(.A(G119), .B(G128), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT24), .B(G110), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(KEYINPUT70), .A3(G110), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n453), .A3(new_n455), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(G119), .B2(new_n204), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n560), .A2(new_n561), .B1(new_n543), .B2(new_n545), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT72), .B(G110), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n552), .A2(new_n553), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n452), .A4(new_n472), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n562), .A2(new_n563), .B1(new_n552), .B2(new_n553), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n452), .A2(new_n472), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT73), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n542), .B1(new_n558), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n568), .A2(new_n571), .ZN(new_n574));
  INV_X1    g388(.A(new_n542), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n557), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n310), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n576), .A3(KEYINPUT25), .A4(new_n310), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n539), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n576), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n574), .B2(new_n557), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n538), .A2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n337), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n335), .A2(G137), .ZN(new_n591));
  OAI21_X1  g405(.A(G131), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n343), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n203), .A2(KEYINPUT65), .A3(new_n205), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT65), .B1(new_n203), .B2(new_n205), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n195), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n344), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(KEYINPUT30), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT30), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n195), .B1(new_n341), .B2(new_n343), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n593), .A2(new_n206), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n262), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n262), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n606), .A3(new_n599), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n458), .A2(G210), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT27), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT26), .B(G101), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT31), .ZN(new_n613));
  INV_X1    g427(.A(new_n611), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT28), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n597), .A2(new_n606), .A3(KEYINPUT28), .A4(new_n599), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n262), .B1(new_n602), .B2(new_n603), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT31), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT66), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT66), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT31), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n310), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT32), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT32), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n626), .A2(new_n630), .A3(new_n627), .A4(new_n310), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT68), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT67), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n593), .B1(new_n365), .B2(new_n366), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n262), .A3(new_n602), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n606), .B1(new_n597), .B2(new_n599), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n634), .B(KEYINPUT28), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n616), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n262), .B1(new_n635), .B2(new_n602), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n607), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n634), .B1(new_n641), .B2(KEYINPUT28), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n611), .A2(KEYINPUT29), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n633), .B1(new_n644), .B2(G902), .ZN(new_n645));
  INV_X1    g459(.A(new_n642), .ZN(new_n646));
  INV_X1    g460(.A(new_n643), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n646), .A2(new_n616), .A3(new_n638), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(KEYINPUT68), .A3(new_n310), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n605), .A2(new_n607), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n614), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT29), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n651), .B(new_n652), .C1(new_n614), .C2(new_n619), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n645), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n589), .B1(new_n632), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n524), .A2(new_n537), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G101), .ZN(G3));
  NOR2_X1   g472(.A1(new_n433), .A2(new_n310), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n432), .B2(new_n433), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n424), .B1(new_n430), .B2(new_n399), .ZN(new_n661));
  INV_X1    g475(.A(new_n399), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n662), .B(new_n425), .C1(new_n429), .C2(new_n419), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT33), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT33), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n426), .A2(new_n431), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(G478), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n515), .A2(new_n521), .ZN(new_n669));
  INV_X1    g483(.A(new_n491), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n314), .A2(new_n313), .A3(new_n324), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n626), .A2(new_n310), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n628), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n589), .A3(new_n533), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT34), .B(G104), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT96), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(new_n488), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n483), .B1(new_n469), .B2(new_n480), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n310), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(KEYINPUT97), .A3(G475), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT97), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n489), .B2(new_n490), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n684), .B(new_n686), .C1(new_n440), .C2(new_n441), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n500), .A2(new_n513), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n689), .A2(new_n516), .B1(new_n514), .B2(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n314), .A2(new_n313), .A3(new_n691), .A4(new_n324), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n676), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NAND2_X1  g509(.A1(new_n579), .A2(new_n580), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n538), .ZN(new_n697));
  OAI22_X1  g511(.A1(new_n558), .A2(new_n572), .B1(KEYINPUT36), .B2(new_n542), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n574), .A2(new_n557), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n585), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT98), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n675), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n524), .A2(new_n537), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  AOI22_X1  g521(.A1(new_n629), .A2(new_n631), .B1(new_n654), .B2(G472), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n697), .A2(new_n702), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n389), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(G900), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n321), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n319), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n687), .A2(new_n690), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n711), .A2(new_n536), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  NOR2_X1   g532(.A1(new_n522), .A2(new_n442), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n314), .A3(new_n703), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n714), .B(KEYINPUT39), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n389), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(KEYINPUT40), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n310), .B1(new_n641), .B2(new_n611), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n650), .A2(new_n611), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n627), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n629), .B2(new_n631), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n313), .B(new_n731), .ZN(new_n732));
  OR3_X1    g546(.A1(new_n725), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G143), .ZN(G45));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n671), .B2(new_n714), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n522), .A2(new_n668), .A3(KEYINPUT100), .A4(new_n715), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n711), .A2(new_n738), .A3(new_n536), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  NOR2_X1   g554(.A1(new_n381), .A2(KEYINPUT101), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n380), .B2(new_n310), .ZN(new_n743));
  AOI211_X1 g557(.A(G902), .B(new_n741), .C1(new_n376), .C2(new_n379), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n329), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n656), .A2(new_n672), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n656), .A2(new_n692), .A3(new_n745), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT102), .B(G116), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G18));
  AND3_X1   g565(.A1(new_n536), .A2(new_n324), .A3(new_n745), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n709), .A2(new_n522), .A3(new_n442), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n632), .B2(new_n655), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  INV_X1    g570(.A(KEYINPUT103), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n697), .A2(new_n757), .A3(new_n586), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT103), .B1(new_n581), .B2(new_n587), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n627), .A2(new_n310), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n621), .B(new_n613), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n614), .B1(new_n639), .B2(new_n642), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n673), .B2(G472), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n760), .A2(new_n719), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n752), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n736), .B2(new_n737), .ZN(new_n770));
  INV_X1    g584(.A(new_n668), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n520), .B(new_n518), .C1(new_n514), .C2(KEYINPUT20), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n771), .B(new_n714), .C1(new_n772), .C2(new_n491), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n671), .A2(new_n735), .A3(new_n714), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(KEYINPUT104), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n536), .A2(new_n745), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n765), .A2(new_n709), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n770), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  INV_X1    g595(.A(new_n760), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n708), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n329), .B1(new_n382), .B2(new_n388), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n314), .A3(new_n312), .A4(new_n303), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n770), .A2(new_n776), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n708), .A2(new_n785), .A3(new_n589), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n776), .A3(new_n770), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n770), .A3(new_n776), .A4(KEYINPUT105), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n786), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n788), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NAND2_X1  g611(.A1(new_n789), .A2(new_n716), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  NAND2_X1  g613(.A1(new_n528), .A2(new_n529), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n387), .A2(KEYINPUT45), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(G469), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT46), .B1(new_n804), .B2(new_n531), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n527), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n531), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n329), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n721), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n772), .A2(new_n491), .A3(new_n668), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT43), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n522), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT43), .B1(new_n814), .B2(new_n668), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n703), .B1(new_n674), .B2(new_n628), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(KEYINPUT44), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n303), .A2(new_n312), .A3(new_n314), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n813), .A2(new_n817), .A3(new_n815), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n810), .A2(new_n818), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G137), .ZN(G39));
  INV_X1    g639(.A(KEYINPUT107), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT47), .B1(new_n808), .B2(new_n809), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n828), .B(new_n329), .C1(new_n806), .C2(new_n807), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n738), .A2(new_n708), .A3(new_n589), .A4(new_n820), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT106), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n827), .A2(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n826), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n827), .A2(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n632), .A2(new_n655), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n588), .A3(new_n819), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(KEYINPUT106), .A3(new_n738), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(KEYINPUT107), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NOR2_X1   g656(.A1(new_n743), .A2(new_n744), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT49), .Z(new_n844));
  NOR4_X1   g658(.A1(new_n844), .A2(new_n535), .A3(new_n330), .A4(new_n782), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n730), .A3(new_n732), .A4(new_n811), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n820), .A2(new_n745), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n588), .A3(new_n320), .A4(new_n730), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n848), .A2(new_n814), .A3(new_n771), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n816), .A2(new_n320), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n779), .A3(new_n847), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n765), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n782), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n743), .A2(new_n744), .A3(new_n526), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n820), .C1(new_n836), .C2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n854), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n732), .A2(new_n535), .A3(new_n745), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n861), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n850), .A3(KEYINPUT50), .A4(new_n854), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT51), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n852), .A3(new_n857), .A4(KEYINPUT51), .ZN(new_n867));
  INV_X1    g681(.A(new_n671), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n316), .B1(new_n848), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n855), .B2(new_n777), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n850), .A2(new_n783), .A3(new_n847), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n785), .A2(new_n778), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n770), .A2(new_n776), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n515), .B1(new_n688), .B2(new_n517), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n686), .A2(new_n684), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n442), .A4(new_n714), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n819), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n837), .A2(new_n883), .A3(new_n389), .A4(new_n709), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT109), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT109), .B1(new_n711), .B2(new_n883), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n798), .B(new_n879), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT108), .B1(new_n814), .B2(new_n442), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT108), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n522), .B(new_n890), .C1(new_n440), .C2(new_n441), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n868), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n676), .A3(new_n536), .A4(new_n324), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n657), .A2(new_n705), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n752), .B1(new_n754), .B2(new_n766), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n746), .A3(new_n749), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n888), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n536), .A2(new_n719), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n709), .A2(new_n715), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n784), .ZN(new_n900));
  INV_X1    g714(.A(new_n729), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n632), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT110), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(new_n900), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n536), .A2(new_n899), .A3(new_n719), .A4(new_n784), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT110), .B1(new_n905), .B2(new_n730), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n711), .B(new_n536), .C1(new_n738), .C2(new_n716), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n780), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT52), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n780), .A3(new_n908), .A4(KEYINPUT52), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n897), .A2(new_n913), .A3(new_n796), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n917));
  XOR2_X1   g731(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n918));
  NAND4_X1  g732(.A1(new_n907), .A2(new_n780), .A3(new_n908), .A4(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n896), .A2(KEYINPUT113), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT113), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n895), .A2(new_n746), .A3(new_n749), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n657), .A2(new_n705), .A3(new_n893), .A4(KEYINPUT53), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n888), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n920), .A2(new_n796), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n916), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n897), .A2(new_n913), .A3(new_n796), .ZN(new_n931));
  INV_X1    g745(.A(new_n915), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n897), .A2(new_n796), .A3(new_n917), .A4(new_n919), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT53), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n877), .B(new_n929), .C1(new_n930), .C2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT116), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n936), .A2(new_n937), .B1(G952), .B2(G953), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n846), .B1(new_n938), .B2(new_n939), .ZN(G75));
  INV_X1    g754(.A(new_n788), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n794), .A2(new_n786), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n792), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n657), .A2(new_n705), .A3(new_n893), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n879), .A2(new_n798), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n895), .A2(new_n746), .A3(new_n749), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n884), .A2(new_n885), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n711), .A2(KEYINPUT109), .A3(new_n883), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n932), .B1(new_n951), .B2(new_n913), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n796), .A2(new_n926), .A3(new_n924), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n917), .A2(new_n919), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(G210), .B(G902), .C1(new_n952), .C2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n271), .A2(new_n278), .A3(new_n213), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n308), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT55), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT117), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(KEYINPUT56), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n956), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n315), .A2(G952), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G51));
  NOR2_X1   g780(.A1(new_n952), .A2(new_n955), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n967), .A2(new_n310), .A3(new_n804), .ZN(new_n968));
  INV_X1    g782(.A(new_n380), .ZN(new_n969));
  INV_X1    g783(.A(new_n928), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n952), .B2(new_n955), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n929), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n383), .B(KEYINPUT57), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT118), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n971), .B2(new_n929), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT118), .B1(new_n978), .B2(new_n969), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n965), .B1(new_n976), .B2(new_n979), .ZN(G54));
  NOR2_X1   g794(.A1(new_n967), .A2(new_n310), .ZN(new_n981));
  NAND2_X1  g795(.A1(KEYINPUT58), .A2(G475), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT119), .Z(new_n983));
  AND3_X1   g797(.A1(new_n981), .A2(new_n689), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n689), .B1(new_n981), .B2(new_n983), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(new_n965), .ZN(G60));
  NAND2_X1  g800(.A1(new_n664), .A2(new_n666), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n659), .B(KEYINPUT59), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n952), .A2(new_n955), .A3(new_n970), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n928), .B1(new_n916), .B2(new_n927), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n965), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n929), .B1(new_n935), .B2(new_n930), .ZN(new_n996));
  INV_X1    g810(.A(new_n989), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT120), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n933), .A2(new_n934), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n951), .A2(new_n932), .A3(new_n913), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n930), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n997), .B1(new_n991), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n988), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT120), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n994), .A4(new_n993), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(new_n1006), .ZN(G63));
  NAND2_X1  g821(.A1(G217), .A2(G902), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT60), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n916), .B2(new_n927), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n698), .A2(new_n700), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n965), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g827(.A1(new_n967), .A2(new_n1009), .B1(new_n582), .B2(new_n583), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT121), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n994), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(KEYINPUT61), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1013), .B(new_n1014), .C1(new_n1017), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(G66));
  OAI21_X1  g836(.A(G953), .B1(new_n322), .B2(new_n210), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n894), .A2(new_n896), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1023), .B1(new_n1024), .B2(G953), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n306), .B(new_n307), .C1(G898), .C2(new_n315), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(G69));
  NAND2_X1  g841(.A1(new_n600), .A2(new_n604), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n492), .A2(new_n493), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT124), .ZN(new_n1031));
  INV_X1    g845(.A(new_n823), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n808), .A2(new_n809), .A3(new_n721), .A4(new_n820), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n821), .A2(new_n822), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n780), .A2(new_n908), .ZN(new_n1036));
  OAI21_X1  g850(.A(KEYINPUT123), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT123), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n824), .A2(new_n1038), .A3(new_n780), .A4(new_n908), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AND2_X1   g854(.A1(new_n810), .A2(new_n898), .ZN(new_n1041));
  AOI22_X1  g855(.A1(new_n1041), .A2(new_n783), .B1(new_n716), .B2(new_n789), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1040), .A2(new_n841), .A3(new_n796), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n315), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n315), .A2(G900), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1031), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g861(.A(KEYINPUT124), .B(new_n1045), .C1(new_n1043), .C2(new_n315), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1030), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(G227), .ZN(new_n1050));
  OAI21_X1  g864(.A(G953), .B1(new_n1050), .B2(new_n712), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n733), .A2(new_n780), .A3(new_n908), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT62), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n722), .A2(new_n819), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n656), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n892), .B(KEYINPUT122), .Z(new_n1057));
  AOI21_X1  g871(.A(new_n1035), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g872(.A1(new_n841), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  OR3_X1    g874(.A1(new_n1060), .A2(G953), .A3(new_n1030), .ZN(new_n1061));
  AND3_X1   g875(.A1(new_n1049), .A2(new_n1051), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1051), .B1(new_n1049), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n1062), .A2(new_n1063), .ZN(G72));
  NOR2_X1   g878(.A1(new_n650), .A2(new_n611), .ZN(new_n1065));
  INV_X1    g879(.A(new_n1024), .ZN(new_n1066));
  OR2_X1    g880(.A1(new_n1043), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT127), .ZN(new_n1068));
  NAND2_X1  g882(.A1(G472), .A2(G902), .ZN(new_n1069));
  XNOR2_X1  g883(.A(new_n1069), .B(KEYINPUT63), .ZN(new_n1070));
  XOR2_X1   g884(.A(new_n1070), .B(KEYINPUT125), .Z(new_n1071));
  AND3_X1   g885(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g886(.A(new_n1068), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1065), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n1054), .A2(new_n1059), .A3(new_n1024), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1075), .A2(new_n1071), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT126), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n1075), .A2(KEYINPUT126), .A3(new_n1071), .ZN(new_n1079));
  NAND4_X1  g893(.A1(new_n1078), .A2(new_n650), .A3(new_n611), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g894(.A(new_n935), .ZN(new_n1081));
  AOI21_X1  g895(.A(new_n1070), .B1(new_n651), .B2(new_n621), .ZN(new_n1082));
  AOI21_X1  g896(.A(new_n965), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g897(.A1(new_n1074), .A2(new_n1080), .A3(new_n1083), .ZN(G57));
endmodule


