//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(G131), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT66), .A2(G137), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT66), .A2(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n193), .A2(KEYINPUT67), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n190), .C1(new_n191), .C2(new_n192), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n189), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT11), .B1(new_n197), .B2(new_n198), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(new_n196), .A3(G137), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n198), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(G137), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT11), .A2(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n203), .A2(new_n210), .A3(G131), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n188), .B1(new_n202), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n193), .A2(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(new_n198), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n201), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT65), .B(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n189), .A3(new_n204), .A4(new_n209), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT70), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n212), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT0), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n222), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n203), .B2(new_n210), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n220), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n228), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT2), .A2(G113), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT2), .A2(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G119), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G116), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G119), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n248), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n241), .A2(new_n243), .B1(new_n245), .B2(new_n220), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n225), .B(new_n231), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n216), .A2(new_n220), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n188), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(new_n221), .ZN(new_n272));
  INV_X1    g086(.A(new_n265), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n248), .A2(new_n265), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n267), .B1(KEYINPUT28), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n279), .B(KEYINPUT27), .Z(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G101), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n228), .B2(new_n247), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n246), .A2(new_n239), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n216), .A2(new_n220), .A3(new_n227), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n289), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n265), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n274), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n289), .A2(new_n290), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n295), .A2(KEYINPUT72), .A3(new_n273), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n272), .A2(new_n297), .A3(new_n273), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n266), .A2(new_n297), .A3(KEYINPUT28), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n294), .B(new_n284), .C1(new_n302), .C2(new_n283), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n187), .B1(new_n286), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n282), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n292), .A2(new_n307), .A3(new_n282), .A4(new_n274), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT32), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  INV_X1    g129(.A(new_n291), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n272), .B2(new_n287), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n266), .B1(new_n317), .B2(new_n265), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n307), .A3(KEYINPUT31), .A4(new_n282), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n308), .A2(new_n309), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n305), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n313), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n314), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n312), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n313), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n304), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n328));
  OR2_X1    g142(.A1(G475), .A2(G902), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n223), .ZN(new_n338));
  OAI211_X1 g152(.A(G146), .B(new_n332), .C1(new_n336), .C2(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G143), .B1(new_n278), .B2(G214), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT17), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT85), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n278), .A2(G214), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n229), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n189), .A3(new_n341), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n341), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT17), .A3(G131), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n338), .A4(new_n339), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n347), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G113), .B(G122), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT18), .A2(G131), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n352), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n362));
  INV_X1    g176(.A(new_n336), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n223), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G146), .B2(new_n336), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n363), .A2(new_n362), .A3(new_n223), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n356), .A2(new_n359), .A3(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT19), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT19), .B1(new_n333), .B2(new_n335), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT84), .B1(new_n371), .B2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n344), .A2(new_n350), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(new_n223), .C1(new_n369), .C2(new_n370), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n372), .A2(new_n339), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n359), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n329), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n328), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n368), .A2(new_n379), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT86), .B1(new_n383), .B2(new_n329), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n259), .A2(G122), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT14), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n388), .B(new_n390), .C1(KEYINPUT14), .C2(new_n386), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n387), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n392));
  OAI21_X1  g206(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n394));
  XNOR2_X1  g208(.A(G128), .B(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n218), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n218), .A2(new_n395), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n390), .A2(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n197), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n396), .A3(KEYINPUT87), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n393), .A2(new_n399), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n400), .B(new_n401), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n229), .A3(G128), .ZN(new_n409));
  OAI211_X1 g223(.A(G134), .B(new_n409), .C1(new_n403), .C2(new_n408), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n410), .A3(new_n396), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT9), .B(G234), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(G953), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT89), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G902), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n422), .B2(new_n423), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT86), .B(new_n328), .C1(new_n383), .C2(new_n329), .ZN(new_n429));
  INV_X1    g243(.A(new_n368), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n359), .B1(new_n356), .B2(new_n367), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G475), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n385), .A2(new_n428), .A3(new_n429), .A4(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(KEYINPUT90), .A2(G952), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT90), .A2(G952), .ZN(new_n437));
  AOI21_X1  g251(.A(G953), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G234), .ZN(new_n439));
  INV_X1    g253(.A(G237), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G953), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n423), .B(new_n442), .C1(G234), .C2(G237), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n434), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G221), .ZN(new_n448));
  INV_X1    g262(.A(new_n412), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n423), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(new_n358), .B2(G107), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n401), .A3(G104), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n358), .A2(G107), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT75), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT75), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n453), .A2(new_n455), .A3(new_n459), .A4(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G101), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G101), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n453), .A2(new_n455), .A3(new_n462), .A4(new_n456), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n452), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n457), .B2(KEYINPUT75), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT4), .B1(new_n465), .B2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n244), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n246), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT76), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n358), .A3(G107), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT76), .B1(new_n358), .B2(G107), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n401), .A2(G104), .ZN(new_n473));
  OAI211_X1 g287(.A(G101), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n269), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n227), .A2(new_n477), .A3(KEYINPUT10), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n467), .A2(new_n468), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n468), .B1(new_n467), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n442), .A2(G227), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n482), .B(new_n483), .Z(new_n484));
  NOR3_X1   g298(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n227), .A2(new_n477), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n269), .A2(new_n475), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n246), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT12), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(KEYINPUT12), .A3(new_n246), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n467), .A2(new_n468), .A3(new_n479), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n486), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n451), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n484), .ZN(new_n499));
  INV_X1    g313(.A(new_n481), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n495), .A3(new_n486), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT77), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n502), .A3(G469), .ZN(new_n503));
  INV_X1    g317(.A(G469), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n423), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n495), .A3(new_n486), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n450), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n447), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g326(.A(G113), .B1(new_n258), .B2(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT78), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n262), .A2(new_n514), .A3(new_n517), .A4(new_n475), .ZN(new_n518));
  XNOR2_X1  g332(.A(G110), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n515), .B1(new_n256), .B2(new_n261), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n475), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n227), .A2(new_n334), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n334), .B2(new_n242), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n442), .A2(G224), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT80), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(KEYINPUT7), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n527), .B2(KEYINPUT7), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n518), .A2(new_n523), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(KEYINPUT7), .A3(new_n526), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n525), .A2(KEYINPUT81), .A3(KEYINPUT7), .A4(new_n526), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n514), .A2(new_n262), .A3(new_n477), .A4(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n461), .A2(new_n463), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n466), .B1(new_n537), .B2(KEYINPUT4), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n536), .B(new_n519), .C1(new_n538), .C2(new_n273), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n538), .B2(new_n273), .ZN(new_n541));
  INV_X1    g355(.A(new_n519), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT6), .A3(new_n539), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n525), .B(new_n526), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n546), .A3(new_n542), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G210), .B1(G237), .B2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT82), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n540), .A2(new_n548), .A3(new_n550), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT82), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n511), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n413), .B1(G234), .B2(new_n423), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n257), .B2(G128), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n566), .A2(KEYINPUT23), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(KEYINPUT23), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n567), .B(new_n568), .C1(G119), .C2(new_n222), .ZN(new_n569));
  XNOR2_X1  g383(.A(G119), .B(G128), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT24), .B(G110), .Z(new_n571));
  OAI22_X1  g385(.A1(new_n569), .A2(G110), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n339), .C1(G146), .C2(new_n336), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n570), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n340), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n448), .A2(new_n439), .A3(G953), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n573), .B2(new_n576), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n564), .B1(new_n584), .B2(G902), .ZN(new_n585));
  OR4_X1    g399(.A1(new_n564), .A2(new_n582), .A3(G902), .A4(new_n583), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n563), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n584), .A2(G902), .A3(new_n562), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n327), .A2(new_n561), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n462), .ZN(G3));
  AOI21_X1  g406(.A(new_n550), .B1(new_n540), .B2(new_n548), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n556), .B1(new_n557), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT92), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n556), .C1(new_n557), .C2(new_n593), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n446), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n429), .A2(new_n433), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n422), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n415), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n424), .A2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n422), .A2(new_n423), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT93), .B(G478), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n385), .A2(new_n600), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n598), .A2(new_n599), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT91), .B(G472), .C1(new_n321), .C2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(KEYINPUT91), .A2(G472), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n312), .A2(new_n423), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n615), .A3(new_n589), .A4(new_n510), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  OAI211_X1 g434(.A(new_n600), .B(new_n385), .C1(new_n427), .C2(new_n426), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n598), .A2(new_n599), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n617), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n577), .B(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n628), .A2(new_n423), .A3(new_n563), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n587), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n511), .A2(new_n559), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n613), .A2(new_n615), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  NAND2_X1  g450(.A1(new_n325), .A2(new_n326), .ZN(new_n637));
  INV_X1    g451(.A(new_n304), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n630), .ZN(new_n640));
  INV_X1    g454(.A(new_n443), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n441), .B1(G900), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT94), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n621), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n598), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n645), .A3(new_n510), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XOR2_X1   g461(.A(new_n643), .B(KEYINPUT39), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n510), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n382), .A2(new_n384), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n429), .A2(new_n433), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n428), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n556), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n555), .A2(new_n558), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT38), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n318), .A2(new_n283), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n423), .B1(new_n276), .B2(new_n282), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n637), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n630), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(new_n606), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n610), .B1(new_n604), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n643), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n667), .B(new_n668), .C1(new_n651), .C2(new_n652), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n595), .A2(new_n670), .A3(new_n597), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT95), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT95), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n595), .A2(new_n670), .A3(new_n673), .A4(new_n597), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n639), .A2(new_n675), .A3(new_n510), .A4(new_n640), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  OR2_X1    g491(.A1(new_n508), .A2(new_n504), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n508), .A2(new_n504), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n450), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT96), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  OR3_X1    g498(.A1(new_n684), .A2(KEYINPUT96), .A3(new_n450), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n639), .A2(new_n612), .A3(new_n589), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n639), .A2(new_n623), .A3(new_n589), .A4(new_n686), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR3_X1   g506(.A1(new_n630), .A2(new_n434), .A3(new_n446), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n684), .A2(new_n450), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n597), .A3(new_n595), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n639), .A2(new_n696), .A3(KEYINPUT98), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n327), .B2(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT99), .B(G119), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n589), .B(new_n703), .ZN(new_n704));
  OAI22_X1  g518(.A1(new_n310), .A2(new_n311), .B1(new_n282), .B2(new_n277), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n313), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n321), .B2(G902), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n598), .A2(new_n654), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n599), .A3(new_n711), .A4(new_n686), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND3_X1  g527(.A1(new_n640), .A2(new_n706), .A3(new_n707), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n671), .A3(new_n682), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n334), .ZN(G27));
  NAND2_X1  g530(.A1(new_n656), .A2(new_n556), .ZN(new_n717));
  INV_X1    g531(.A(new_n679), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n505), .B(KEYINPUT101), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n499), .A2(new_n501), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n720), .B2(new_n504), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n681), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n669), .A2(KEYINPUT42), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n639), .A2(new_n589), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n670), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n638), .A2(new_n314), .A3(new_n323), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n704), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT102), .B(G131), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G33));
  NAND4_X1  g546(.A1(new_n639), .A2(new_n589), .A3(new_n644), .A4(new_n723), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND2_X1  g548(.A1(new_n632), .A2(new_n640), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n632), .A2(KEYINPUT105), .A3(new_n640), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n653), .A2(new_n667), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n556), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n555), .B2(new_n558), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n739), .A2(KEYINPUT44), .A3(new_n742), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n751), .A3(new_n748), .A4(new_n747), .ZN(new_n752));
  INV_X1    g566(.A(new_n719), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n497), .A2(new_n502), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n720), .B2(new_n755), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT103), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n497), .B2(new_n502), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT103), .B1(new_n761), .B2(new_n757), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n753), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n718), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n719), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n764), .A2(KEYINPUT104), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n679), .B1(new_n767), .B2(new_n765), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n450), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n750), .A2(new_n648), .A3(new_n752), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  XNOR2_X1  g588(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n772), .B(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n639), .A2(new_n589), .A3(new_n669), .A4(new_n717), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n768), .A2(new_n771), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n781), .B2(new_n450), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n775), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  NAND3_X1  g601(.A1(new_n704), .A2(new_n556), .A3(new_n681), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n684), .B(KEYINPUT49), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n740), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n663), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n657), .ZN(new_n792));
  INV_X1    g606(.A(new_n714), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n723), .A3(new_n670), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n510), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n327), .A2(new_n796), .A3(new_n630), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n434), .A2(KEYINPUT110), .A3(new_n643), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT110), .B1(new_n434), .B2(new_n643), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n798), .A2(new_n747), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n795), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n730), .A2(new_n733), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n700), .A2(new_n687), .A3(new_n691), .A4(new_n712), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n560), .A2(new_n640), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n600), .A2(new_n385), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n667), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n446), .B1(new_n806), .B2(new_n621), .ZN(new_n807));
  INV_X1    g621(.A(new_n559), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n804), .A2(new_n632), .B1(new_n616), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT109), .B1(new_n591), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n639), .A2(new_n589), .A3(new_n560), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n813));
  INV_X1    g627(.A(new_n809), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n814), .A2(new_n617), .B1(new_n631), .B2(new_n633), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n802), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n722), .A2(new_n643), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n597), .A2(new_n819), .A3(new_n595), .A4(new_n654), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n663), .A2(new_n630), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n715), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n676), .A2(new_n646), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n327), .A2(new_n796), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n715), .B1(new_n825), .B2(new_n645), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n676), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n818), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT98), .B1(new_n639), .B2(new_n696), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n327), .A2(new_n695), .A3(new_n698), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n691), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n712), .A2(new_n687), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n591), .A2(new_n810), .A3(KEYINPUT109), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n725), .A2(new_n733), .A3(new_n729), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n639), .A2(new_n800), .A3(new_n510), .A4(new_n640), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n794), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n829), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n831), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n818), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n844), .B2(new_n829), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT111), .A4(new_n851), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n441), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n742), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT112), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n717), .A2(new_n682), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n793), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n791), .A2(new_n589), .A3(new_n856), .A4(new_n859), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n653), .A2(new_n610), .A3(new_n607), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n710), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n657), .A2(new_n746), .A3(new_n694), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n866), .A2(KEYINPUT50), .A3(new_n868), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n747), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT113), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n777), .B1(new_n450), .B2(new_n680), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n438), .B(KEYINPUT116), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n598), .A2(new_n694), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n860), .A2(new_n704), .A3(new_n727), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n887));
  OAI221_X1 g701(.A(new_n884), .B1(new_n885), .B2(new_n865), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n806), .B2(new_n862), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n855), .A2(new_n882), .A3(new_n883), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n792), .B1(new_n891), .B2(new_n892), .ZN(G75));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n849), .A2(new_n850), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G902), .ZN(new_n896));
  INV_X1    g710(.A(G210), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n544), .A2(new_n547), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(new_n545), .Z(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n901), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n442), .A2(G952), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT118), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT119), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(G51));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n847), .A2(new_n908), .A3(new_n852), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n895), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n719), .B(KEYINPUT57), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n506), .A2(new_n507), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n896), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n766), .B(KEYINPUT121), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n914), .B2(new_n917), .ZN(G54));
  INV_X1    g732(.A(new_n383), .ZN(new_n919));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n896), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n896), .B2(new_n920), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n905), .B1(new_n921), .B2(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n853), .A2(new_n854), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n604), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n909), .A2(new_n605), .A3(new_n910), .A4(new_n926), .ZN(new_n929));
  INV_X1    g743(.A(new_n906), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n604), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n934), .A3(new_n930), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n895), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n584), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n895), .A2(new_n628), .A3(new_n939), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n930), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT61), .Z(G66));
  INV_X1    g758(.A(G224), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n444), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n803), .A2(new_n817), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n899), .B1(G898), .B2(new_n442), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n317), .B(new_n371), .Z(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(G900), .B2(new_n442), .ZN(new_n953));
  INV_X1    g767(.A(new_n728), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n772), .A2(new_n648), .A3(new_n711), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n676), .A3(new_n826), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n840), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n786), .A2(new_n773), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n953), .B1(new_n958), .B2(new_n442), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n952), .A2(G953), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n649), .B(new_n717), .C1(new_n806), .C2(new_n621), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n639), .A3(new_n589), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n773), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n664), .A2(new_n826), .A3(new_n676), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n780), .A2(new_n785), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n960), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n951), .B1(new_n959), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n951), .C1(new_n959), .C2(new_n969), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n442), .B1(G227), .B2(G900), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n971), .B2(new_n973), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  NAND4_X1  g791(.A1(new_n786), .A2(new_n773), .A3(new_n947), .A4(new_n957), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n187), .A2(new_n423), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(new_n981));
  AOI211_X1 g795(.A(new_n282), .B(new_n293), .C1(new_n978), .C2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT127), .B1(new_n982), .B2(new_n905), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n963), .A2(new_n968), .A3(new_n947), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n981), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n318), .A2(new_n282), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n294), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n985), .A2(new_n660), .B1(new_n895), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n905), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G57));
endmodule


