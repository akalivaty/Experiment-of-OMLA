

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  INV_X1 U373 ( .A(n644), .ZN(n351) );
  AND2_X1 U374 ( .A1(n718), .A2(G472), .ZN(n641) );
  NAND2_X1 U375 ( .A1(n602), .A2(n601), .ZN(n432) );
  XNOR2_X1 U376 ( .A(n526), .B(n525), .ZN(n569) );
  XNOR2_X1 U377 ( .A(n353), .B(n410), .ZN(n713) );
  XNOR2_X1 U378 ( .A(n737), .B(n520), .ZN(n353) );
  XNOR2_X1 U379 ( .A(n377), .B(n521), .ZN(n737) );
  XNOR2_X1 U380 ( .A(n352), .B(n351), .ZN(G57) );
  NAND2_X1 U381 ( .A1(n428), .A2(n427), .ZN(n352) );
  XNOR2_X2 U382 ( .A(n570), .B(KEYINPUT19), .ZN(n602) );
  XNOR2_X2 U383 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n376) );
  NOR2_X1 U384 ( .A1(G237), .A2(G953), .ZN(n479) );
  OR2_X1 U385 ( .A1(n454), .A2(n453), .ZN(n660) );
  XNOR2_X2 U386 ( .A(n495), .B(n494), .ZN(n614) );
  NOR2_X2 U387 ( .A1(n625), .A2(n435), .ZN(n605) );
  AND2_X1 U388 ( .A1(n417), .A2(n363), .ZN(n415) );
  NOR2_X1 U389 ( .A1(n757), .A2(KEYINPUT44), .ZN(n423) );
  AND2_X1 U390 ( .A1(n576), .A2(n692), .ZN(n528) );
  AND2_X1 U391 ( .A1(n513), .A2(n512), .ZN(n576) );
  AND2_X1 U392 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U393 ( .A(n554), .B(n457), .ZN(n663) );
  NAND2_X1 U394 ( .A1(n395), .A2(n393), .ZN(n406) );
  XNOR2_X1 U395 ( .A(n739), .B(n471), .ZN(n514) );
  XNOR2_X1 U396 ( .A(n503), .B(n502), .ZN(n739) );
  NAND2_X1 U397 ( .A1(n713), .A2(n710), .ZN(n526) );
  XNOR2_X1 U398 ( .A(n437), .B(n436), .ZN(n619) );
  AND2_X1 U399 ( .A1(n402), .A2(n399), .ZN(n631) );
  XNOR2_X2 U400 ( .A(n432), .B(n603), .ZN(n623) );
  NOR2_X1 U401 ( .A1(n582), .A2(n581), .ZN(n588) );
  INV_X1 U402 ( .A(n672), .ZN(n462) );
  XNOR2_X1 U403 ( .A(n543), .B(n359), .ZN(n748) );
  NAND2_X1 U404 ( .A1(n391), .A2(n433), .ZN(n622) );
  INV_X1 U405 ( .A(G472), .ZN(n385) );
  OR2_X1 U406 ( .A1(n642), .A2(G902), .ZN(n386) );
  XNOR2_X1 U407 ( .A(n538), .B(n440), .ZN(n722) );
  XNOR2_X1 U408 ( .A(n539), .B(n540), .ZN(n440) );
  INV_X1 U409 ( .A(n514), .ZN(n398) );
  XNOR2_X1 U410 ( .A(KEYINPUT15), .B(G902), .ZN(n710) );
  AND2_X1 U411 ( .A1(n638), .A2(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U412 ( .A(n636), .B(n461), .ZN(n638) );
  XNOR2_X1 U413 ( .A(n613), .B(n365), .ZN(n402) );
  NAND2_X1 U414 ( .A1(n406), .A2(n405), .ZN(n404) );
  NOR2_X1 U415 ( .A1(n355), .A2(G902), .ZN(n405) );
  INV_X1 U416 ( .A(KEYINPUT92), .ZN(n436) );
  NOR2_X2 U417 ( .A1(n758), .A2(n653), .ZN(n437) );
  XOR2_X1 U418 ( .A(KEYINPUT104), .B(KEYINPUT11), .Z(n533) );
  XNOR2_X1 U419 ( .A(G122), .B(G140), .ZN(n532) );
  XOR2_X1 U420 ( .A(G113), .B(G104), .Z(n531) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(G137), .Z(n476) );
  INV_X1 U422 ( .A(G140), .ZN(n375) );
  XOR2_X1 U423 ( .A(KEYINPUT9), .B(G122), .Z(n545) );
  OR2_X2 U424 ( .A1(n473), .A2(G134), .ZN(n474) );
  XNOR2_X1 U425 ( .A(G116), .B(G113), .ZN(n478) );
  XOR2_X1 U426 ( .A(G119), .B(KEYINPUT3), .Z(n360) );
  INV_X1 U427 ( .A(KEYINPUT109), .ZN(n455) );
  NOR2_X1 U428 ( .A1(n663), .A2(n665), .ZN(n456) );
  NAND2_X1 U429 ( .A1(n414), .A2(n413), .ZN(n636) );
  NAND2_X1 U430 ( .A1(n418), .A2(n419), .ZN(n413) );
  AND2_X1 U431 ( .A1(n416), .A2(n415), .ZN(n414) );
  NAND2_X1 U432 ( .A1(n692), .A2(n691), .ZN(n412) );
  XNOR2_X1 U433 ( .A(n524), .B(KEYINPUT95), .ZN(n525) );
  INV_X1 U434 ( .A(KEYINPUT1), .ZN(n392) );
  AND2_X1 U435 ( .A1(n584), .A2(n381), .ZN(n380) );
  INV_X1 U436 ( .A(KEYINPUT83), .ZN(n384) );
  INV_X1 U437 ( .A(KEYINPUT0), .ZN(n603) );
  NAND2_X1 U438 ( .A1(n569), .A2(n691), .ZN(n570) );
  XNOR2_X1 U439 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U440 ( .A(KEYINPUT25), .ZN(n492) );
  XNOR2_X1 U441 ( .A(n541), .B(n439), .ZN(n558) );
  XNOR2_X1 U442 ( .A(n542), .B(G475), .ZN(n439) );
  NAND2_X1 U443 ( .A1(n718), .A2(n468), .ZN(n469) );
  AND2_X1 U444 ( .A1(n711), .A2(n372), .ZN(n468) );
  XOR2_X1 U445 ( .A(n552), .B(n551), .Z(n723) );
  XNOR2_X1 U446 ( .A(n398), .B(n463), .ZN(n394) );
  INV_X1 U447 ( .A(G953), .ZN(n750) );
  XNOR2_X1 U448 ( .A(n568), .B(n567), .ZN(n420) );
  OR2_X1 U449 ( .A1(G902), .A2(G237), .ZN(n523) );
  XNOR2_X1 U450 ( .A(n490), .B(n434), .ZN(n496) );
  XNOR2_X1 U451 ( .A(n491), .B(KEYINPUT100), .ZN(n434) );
  XOR2_X1 U452 ( .A(KEYINPUT101), .B(KEYINPUT20), .Z(n491) );
  INV_X1 U453 ( .A(KEYINPUT73), .ZN(n421) );
  XNOR2_X1 U454 ( .A(n517), .B(KEYINPUT10), .ZN(n536) );
  XNOR2_X1 U455 ( .A(G143), .B(G131), .ZN(n530) );
  NAND2_X1 U456 ( .A1(G237), .A2(G234), .ZN(n506) );
  AND2_X1 U457 ( .A1(n680), .A2(n357), .ZN(n459) );
  XNOR2_X1 U458 ( .A(n449), .B(KEYINPUT69), .ZN(n584) );
  NAND2_X1 U459 ( .A1(n614), .A2(n450), .ZN(n449) );
  AND2_X1 U460 ( .A1(n560), .A2(n357), .ZN(n450) );
  NAND2_X1 U461 ( .A1(n355), .A2(G902), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n356), .B(n477), .ZN(n441) );
  XNOR2_X1 U463 ( .A(G110), .B(G107), .ZN(n503) );
  XNOR2_X1 U464 ( .A(n447), .B(n446), .ZN(n484) );
  XNOR2_X1 U465 ( .A(G119), .B(KEYINPUT80), .ZN(n446) );
  XNOR2_X1 U466 ( .A(n448), .B(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U467 ( .A(KEYINPUT99), .B(KEYINPUT24), .ZN(n448) );
  XOR2_X1 U468 ( .A(n536), .B(n500), .Z(n747) );
  XNOR2_X1 U469 ( .A(n636), .B(n445), .ZN(n749) );
  INV_X1 U470 ( .A(KEYINPUT85), .ZN(n445) );
  XNOR2_X1 U471 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n486) );
  XNOR2_X1 U472 ( .A(G107), .B(G116), .ZN(n544) );
  XNOR2_X1 U473 ( .A(n501), .B(n499), .ZN(n463) );
  XNOR2_X1 U474 ( .A(n362), .B(n398), .ZN(n396) );
  XNOR2_X1 U475 ( .A(n748), .B(G146), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n515), .B(n516), .ZN(n470) );
  XNOR2_X1 U477 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n516) );
  XNOR2_X1 U478 ( .A(n376), .B(G122), .ZN(n522) );
  XNOR2_X1 U479 ( .A(n442), .B(n366), .ZN(n435) );
  NOR2_X1 U480 ( .A1(n622), .A2(n630), .ZN(n442) );
  INV_X1 U481 ( .A(n399), .ZN(n391) );
  NOR2_X1 U482 ( .A1(n412), .A2(n694), .ZN(n559) );
  INV_X1 U483 ( .A(KEYINPUT98), .ZN(n604) );
  BUF_X1 U484 ( .A(n680), .Z(n433) );
  AND2_X1 U485 ( .A1(n711), .A2(n371), .ZN(n464) );
  XNOR2_X1 U486 ( .A(n514), .B(n411), .ZN(n410) );
  XNOR2_X1 U487 ( .A(n470), .B(KEYINPUT81), .ZN(n411) );
  NOR2_X1 U488 ( .A1(n593), .A2(n590), .ZN(n585) );
  INV_X1 U489 ( .A(KEYINPUT32), .ZN(n400) );
  NAND2_X1 U490 ( .A1(n458), .A2(n438), .ZN(n453) );
  BUF_X1 U491 ( .A(n602), .Z(n438) );
  NOR2_X1 U492 ( .A1(n628), .A2(n467), .ZN(n466) );
  INV_X1 U493 ( .A(KEYINPUT108), .ZN(n457) );
  NOR2_X1 U494 ( .A1(n678), .A2(n632), .ZN(n646) );
  XNOR2_X1 U495 ( .A(n379), .B(n378), .ZN(n632) );
  INV_X1 U496 ( .A(KEYINPUT89), .ZN(n378) );
  INV_X1 U497 ( .A(KEYINPUT121), .ZN(n425) );
  XNOR2_X1 U498 ( .A(n469), .B(n723), .ZN(n724) );
  INV_X1 U499 ( .A(KEYINPUT60), .ZN(n429) );
  XNOR2_X1 U500 ( .A(n720), .B(n443), .ZN(n721) );
  XOR2_X1 U501 ( .A(n505), .B(G469), .Z(n355) );
  XNOR2_X1 U502 ( .A(n375), .B(G137), .ZN(n500) );
  XOR2_X1 U503 ( .A(n521), .B(n480), .Z(n356) );
  OR2_X1 U504 ( .A1(n598), .A2(n511), .ZN(n357) );
  AND2_X1 U505 ( .A1(n621), .A2(n388), .ZN(n358) );
  XOR2_X1 U506 ( .A(G131), .B(KEYINPUT4), .Z(n359) );
  AND2_X1 U507 ( .A1(n663), .A2(n380), .ZN(n361) );
  XOR2_X1 U508 ( .A(n501), .B(n499), .Z(n362) );
  INV_X1 U509 ( .A(n564), .ZN(n458) );
  AND2_X1 U510 ( .A1(n673), .A2(n462), .ZN(n363) );
  XNOR2_X1 U511 ( .A(n562), .B(n561), .ZN(n364) );
  XOR2_X1 U512 ( .A(n612), .B(KEYINPUT22), .Z(n365) );
  XOR2_X1 U513 ( .A(n596), .B(n595), .Z(n366) );
  XNOR2_X1 U514 ( .A(KEYINPUT48), .B(KEYINPUT68), .ZN(n367) );
  XOR2_X1 U515 ( .A(n642), .B(KEYINPUT62), .Z(n368) );
  XNOR2_X1 U516 ( .A(n722), .B(KEYINPUT59), .ZN(n369) );
  NOR2_X1 U517 ( .A1(n710), .A2(n709), .ZN(n370) );
  AND2_X1 U518 ( .A1(n640), .A2(G217), .ZN(n371) );
  AND2_X1 U519 ( .A1(n640), .A2(G478), .ZN(n372) );
  XNOR2_X1 U520 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n373) );
  INV_X1 U521 ( .A(KEYINPUT86), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n426), .B(n425), .ZN(G63) );
  NOR2_X1 U523 ( .A1(n614), .A2(n610), .ZN(n680) );
  NOR2_X1 U524 ( .A1(n729), .A2(n728), .ZN(n730) );
  INV_X1 U525 ( .A(n728), .ZN(n427) );
  NOR2_X1 U526 ( .A1(n724), .A2(n728), .ZN(n426) );
  NAND2_X1 U527 ( .A1(n374), .A2(n355), .ZN(n409) );
  INV_X1 U528 ( .A(n406), .ZN(n374) );
  XNOR2_X1 U529 ( .A(n406), .B(n373), .ZN(n443) );
  XNOR2_X2 U530 ( .A(n360), .B(n478), .ZN(n521) );
  XNOR2_X1 U531 ( .A(n522), .B(KEYINPUT16), .ZN(n377) );
  AND2_X2 U532 ( .A1(n631), .A2(n466), .ZN(n653) );
  NAND2_X1 U533 ( .A1(n631), .A2(n630), .ZN(n379) );
  AND2_X1 U534 ( .A1(n634), .A2(n620), .ZN(n388) );
  INV_X1 U535 ( .A(n473), .ZN(n515) );
  INV_X1 U536 ( .A(n630), .ZN(n381) );
  INV_X1 U537 ( .A(n587), .ZN(n669) );
  OR2_X1 U538 ( .A1(n586), .A2(n616), .ZN(n587) );
  NAND2_X2 U539 ( .A1(n407), .A2(n404), .ZN(n583) );
  NAND2_X1 U540 ( .A1(n403), .A2(n394), .ZN(n393) );
  XNOR2_X2 U541 ( .A(n382), .B(n421), .ZN(n389) );
  NAND2_X1 U542 ( .A1(n424), .A2(n422), .ZN(n382) );
  NAND2_X1 U543 ( .A1(n402), .A2(n383), .ZN(n401) );
  XNOR2_X1 U544 ( .A(n617), .B(n384), .ZN(n383) );
  XNOR2_X2 U545 ( .A(n386), .B(n385), .ZN(n683) );
  XNOR2_X2 U546 ( .A(n387), .B(KEYINPUT45), .ZN(n734) );
  NAND2_X2 U547 ( .A1(n389), .A2(n358), .ZN(n387) );
  XNOR2_X2 U548 ( .A(G143), .B(G128), .ZN(n473) );
  AND2_X1 U549 ( .A1(n390), .A2(n399), .ZN(n681) );
  INV_X1 U550 ( .A(n433), .ZN(n390) );
  XNOR2_X1 U551 ( .A(n399), .B(KEYINPUT94), .ZN(n616) );
  NOR2_X1 U552 ( .A1(n590), .A2(n391), .ZN(n592) );
  XNOR2_X2 U553 ( .A(n583), .B(n392), .ZN(n399) );
  NAND2_X1 U554 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U555 ( .A(n403), .ZN(n397) );
  XNOR2_X2 U556 ( .A(n401), .B(n400), .ZN(n758) );
  XNOR2_X1 U557 ( .A(n441), .B(n403), .ZN(n642) );
  NOR2_X1 U558 ( .A1(n695), .A2(n412), .ZN(n696) );
  NAND2_X1 U559 ( .A1(n420), .A2(n367), .ZN(n416) );
  NAND2_X1 U560 ( .A1(n589), .A2(n367), .ZN(n417) );
  NOR2_X1 U561 ( .A1(n589), .A2(n367), .ZN(n418) );
  INV_X1 U562 ( .A(n420), .ZN(n419) );
  XNOR2_X1 U563 ( .A(n423), .B(KEYINPUT66), .ZN(n422) );
  XNOR2_X1 U564 ( .A(n619), .B(KEYINPUT91), .ZN(n424) );
  NAND2_X1 U565 ( .A1(n725), .A2(G475), .ZN(n444) );
  NAND2_X2 U566 ( .A1(n465), .A2(n637), .ZN(n718) );
  XNOR2_X1 U567 ( .A(n643), .B(n368), .ZN(n428) );
  XNOR2_X1 U568 ( .A(n430), .B(n429), .ZN(G60) );
  NAND2_X1 U569 ( .A1(n431), .A2(n427), .ZN(n430) );
  XNOR2_X1 U570 ( .A(n444), .B(n369), .ZN(n431) );
  AND2_X2 U571 ( .A1(n719), .A2(n718), .ZN(n725) );
  XNOR2_X1 U572 ( .A(n460), .B(KEYINPUT79), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n489), .B(n488), .ZN(n727) );
  NOR2_X1 U574 ( .A1(n555), .A2(n661), .ZN(n557) );
  NAND2_X1 U575 ( .A1(n623), .A2(n611), .ZN(n613) );
  INV_X1 U576 ( .A(n695), .ZN(n451) );
  XOR2_X2 U577 ( .A(n683), .B(KEYINPUT6), .Z(n630) );
  NOR2_X1 U578 ( .A1(G902), .A2(n727), .ZN(n495) );
  NOR2_X1 U579 ( .A1(n749), .A2(n461), .ZN(n635) );
  NAND2_X2 U580 ( .A1(n474), .A2(n475), .ZN(n543) );
  INV_X1 U581 ( .A(n504), .ZN(n471) );
  AND2_X2 U582 ( .A1(n711), .A2(n640), .ZN(n719) );
  XNOR2_X1 U583 ( .A(n563), .B(n364), .ZN(n454) );
  INV_X1 U584 ( .A(n660), .ZN(n452) );
  NAND2_X1 U585 ( .A1(n452), .A2(n451), .ZN(n572) );
  XNOR2_X2 U586 ( .A(n456), .B(n455), .ZN(n695) );
  NOR2_X1 U587 ( .A1(n454), .A2(n564), .ZN(n571) );
  NAND2_X1 U588 ( .A1(n459), .A2(n583), .ZN(n460) );
  NAND2_X1 U589 ( .A1(n583), .A2(n433), .ZN(n626) );
  NAND2_X1 U590 ( .A1(n718), .A2(n464), .ZN(n726) );
  NAND2_X1 U591 ( .A1(n635), .A2(n734), .ZN(n465) );
  INV_X1 U592 ( .A(n614), .ZN(n467) );
  NAND2_X2 U593 ( .A1(n734), .A2(n639), .ZN(n711) );
  XNOR2_X1 U594 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n472) );
  INV_X1 U595 ( .A(KEYINPUT93), .ZN(n595) );
  INV_X1 U596 ( .A(G104), .ZN(n502) );
  INV_X1 U597 ( .A(KEYINPUT28), .ZN(n561) );
  XNOR2_X1 U598 ( .A(n713), .B(n472), .ZN(n714) );
  XNOR2_X1 U599 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U600 ( .A1(G952), .A2(n750), .ZN(n728) );
  INV_X1 U601 ( .A(KEYINPUT30), .ZN(n482) );
  NAND2_X1 U602 ( .A1(n473), .A2(G134), .ZN(n475) );
  XOR2_X1 U603 ( .A(KEYINPUT65), .B(G101), .Z(n504) );
  XNOR2_X1 U604 ( .A(n476), .B(n504), .ZN(n477) );
  XNOR2_X1 U605 ( .A(n479), .B(KEYINPUT78), .ZN(n529) );
  NAND2_X1 U606 ( .A1(G210), .A2(n529), .ZN(n480) );
  INV_X1 U607 ( .A(n683), .ZN(n628) );
  NAND2_X1 U608 ( .A1(G214), .A2(n523), .ZN(n691) );
  NAND2_X1 U609 ( .A1(n628), .A2(n691), .ZN(n481) );
  XNOR2_X1 U610 ( .A(n482), .B(n481), .ZN(n513) );
  XNOR2_X2 U611 ( .A(G125), .B(G146), .ZN(n517) );
  XNOR2_X1 U612 ( .A(G128), .B(G110), .ZN(n483) );
  XNOR2_X1 U613 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U614 ( .A(n747), .B(n485), .ZN(n489) );
  NAND2_X1 U615 ( .A1(n750), .A2(G234), .ZN(n487) );
  XNOR2_X1 U616 ( .A(n487), .B(n486), .ZN(n548) );
  AND2_X1 U617 ( .A1(G221), .A2(n548), .ZN(n488) );
  NAND2_X1 U618 ( .A1(G234), .A2(n710), .ZN(n490) );
  NAND2_X1 U619 ( .A1(G217), .A2(n496), .ZN(n493) );
  XOR2_X1 U620 ( .A(KEYINPUT102), .B(KEYINPUT21), .Z(n498) );
  NAND2_X1 U621 ( .A1(G221), .A2(n496), .ZN(n497) );
  XOR2_X1 U622 ( .A(n498), .B(n497), .Z(n677) );
  XOR2_X1 U623 ( .A(n677), .B(KEYINPUT103), .Z(n610) );
  INV_X1 U624 ( .A(n500), .ZN(n499) );
  NAND2_X1 U625 ( .A1(G227), .A2(n750), .ZN(n501) );
  XNOR2_X1 U626 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n505) );
  XNOR2_X1 U627 ( .A(n506), .B(KEYINPUT96), .ZN(n507) );
  XNOR2_X1 U628 ( .A(KEYINPUT14), .B(n507), .ZN(n508) );
  NAND2_X1 U629 ( .A1(G952), .A2(n508), .ZN(n703) );
  NOR2_X1 U630 ( .A1(G953), .A2(n703), .ZN(n598) );
  NAND2_X1 U631 ( .A1(n508), .A2(G902), .ZN(n509) );
  XNOR2_X1 U632 ( .A(n509), .B(KEYINPUT97), .ZN(n597) );
  NAND2_X1 U633 ( .A1(G953), .A2(n597), .ZN(n510) );
  NOR2_X1 U634 ( .A1(G900), .A2(n510), .ZN(n511) );
  XNOR2_X1 U635 ( .A(n517), .B(KEYINPUT18), .ZN(n519) );
  NAND2_X1 U636 ( .A1(G224), .A2(n750), .ZN(n518) );
  XOR2_X1 U637 ( .A(n519), .B(n518), .Z(n520) );
  NAND2_X1 U638 ( .A1(n523), .A2(G210), .ZN(n524) );
  INV_X1 U639 ( .A(n569), .ZN(n593) );
  XNOR2_X1 U640 ( .A(n593), .B(KEYINPUT38), .ZN(n692) );
  XNOR2_X1 U641 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n527) );
  XNOR2_X1 U642 ( .A(n528), .B(n527), .ZN(n555) );
  XNOR2_X1 U643 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n542) );
  NAND2_X1 U644 ( .A1(n529), .A2(G214), .ZN(n540) );
  XNOR2_X1 U645 ( .A(n531), .B(n530), .ZN(n535) );
  XNOR2_X1 U646 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U647 ( .A(n535), .B(n534), .ZN(n539) );
  XNOR2_X1 U648 ( .A(n536), .B(KEYINPUT12), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n537), .B(KEYINPUT105), .ZN(n538) );
  NOR2_X1 U650 ( .A1(G902), .A2(n722), .ZN(n541) );
  XNOR2_X1 U651 ( .A(KEYINPUT107), .B(KEYINPUT7), .ZN(n552) );
  INV_X1 U652 ( .A(n543), .ZN(n547) );
  XNOR2_X1 U653 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n547), .B(n546), .ZN(n550) );
  NAND2_X1 U655 ( .A1(G217), .A2(n548), .ZN(n549) );
  XNOR2_X1 U656 ( .A(n550), .B(n549), .ZN(n551) );
  NOR2_X1 U657 ( .A1(G902), .A2(n723), .ZN(n553) );
  XNOR2_X1 U658 ( .A(G478), .B(n553), .ZN(n574) );
  NOR2_X1 U659 ( .A1(n558), .A2(n574), .ZN(n665) );
  INV_X1 U660 ( .A(n665), .ZN(n654) );
  NOR2_X1 U661 ( .A1(n555), .A2(n654), .ZN(n672) );
  NAND2_X1 U662 ( .A1(n558), .A2(n574), .ZN(n554) );
  INV_X1 U663 ( .A(n663), .ZN(n661) );
  INV_X1 U664 ( .A(KEYINPUT40), .ZN(n556) );
  XNOR2_X1 U665 ( .A(n557), .B(n556), .ZN(n761) );
  INV_X1 U666 ( .A(n558), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n573), .A2(n574), .ZN(n694) );
  XNOR2_X1 U668 ( .A(KEYINPUT41), .B(n559), .ZN(n690) );
  INV_X1 U669 ( .A(n690), .ZN(n565) );
  INV_X1 U670 ( .A(n677), .ZN(n560) );
  AND2_X1 U671 ( .A1(n584), .A2(n628), .ZN(n563) );
  INV_X1 U672 ( .A(KEYINPUT113), .ZN(n562) );
  XOR2_X1 U673 ( .A(n583), .B(KEYINPUT112), .Z(n564) );
  NAND2_X1 U674 ( .A1(n565), .A2(n571), .ZN(n566) );
  XNOR2_X1 U675 ( .A(KEYINPUT42), .B(n566), .ZN(n759) );
  NAND2_X1 U676 ( .A1(n761), .A2(n759), .ZN(n568) );
  XOR2_X1 U677 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n567) );
  NAND2_X1 U678 ( .A1(n572), .A2(KEYINPUT47), .ZN(n577) );
  OR2_X1 U679 ( .A1(n574), .A2(n573), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n593), .A2(n606), .ZN(n575) );
  NAND2_X1 U681 ( .A1(n576), .A2(n575), .ZN(n659) );
  NAND2_X1 U682 ( .A1(n577), .A2(n659), .ZN(n578) );
  XNOR2_X1 U683 ( .A(n578), .B(KEYINPUT84), .ZN(n582) );
  NOR2_X1 U684 ( .A1(n695), .A2(KEYINPUT47), .ZN(n579) );
  XNOR2_X1 U685 ( .A(KEYINPUT77), .B(n579), .ZN(n580) );
  NOR2_X1 U686 ( .A1(n660), .A2(n580), .ZN(n581) );
  NAND2_X1 U687 ( .A1(n361), .A2(n691), .ZN(n590) );
  XOR2_X1 U688 ( .A(KEYINPUT36), .B(n585), .Z(n586) );
  NAND2_X1 U689 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U690 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n591) );
  XNOR2_X1 U691 ( .A(n592), .B(n591), .ZN(n594) );
  NAND2_X1 U692 ( .A1(n594), .A2(n593), .ZN(n673) );
  XOR2_X1 U693 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n596) );
  NOR2_X1 U694 ( .A1(G898), .A2(n750), .ZN(n742) );
  NAND2_X1 U695 ( .A1(n742), .A2(n597), .ZN(n600) );
  INV_X1 U696 ( .A(n598), .ZN(n599) );
  NAND2_X1 U697 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U698 ( .A(n623), .B(n604), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n605), .B(KEYINPUT34), .ZN(n608) );
  XOR2_X1 U700 ( .A(KEYINPUT82), .B(n606), .Z(n607) );
  NAND2_X1 U701 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X2 U702 ( .A(n609), .B(KEYINPUT35), .ZN(n757) );
  NOR2_X1 U703 ( .A1(n610), .A2(n694), .ZN(n611) );
  XNOR2_X1 U704 ( .A(KEYINPUT64), .B(KEYINPUT74), .ZN(n612) );
  XNOR2_X1 U705 ( .A(n614), .B(KEYINPUT110), .ZN(n678) );
  NAND2_X1 U706 ( .A1(n630), .A2(n678), .ZN(n615) );
  NOR2_X1 U707 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U708 ( .A1(n757), .A2(KEYINPUT44), .ZN(n618) );
  XNOR2_X1 U709 ( .A(n618), .B(KEYINPUT90), .ZN(n621) );
  NAND2_X1 U710 ( .A1(n619), .A2(KEYINPUT44), .ZN(n620) );
  NOR2_X1 U711 ( .A1(n683), .A2(n622), .ZN(n687) );
  NAND2_X1 U712 ( .A1(n623), .A2(n687), .ZN(n624) );
  XNOR2_X1 U713 ( .A(n624), .B(KEYINPUT31), .ZN(n666) );
  OR2_X1 U714 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U715 ( .A1(n628), .A2(n627), .ZN(n648) );
  NOR2_X1 U716 ( .A1(n666), .A2(n648), .ZN(n629) );
  NOR2_X1 U717 ( .A1(n695), .A2(n629), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n633), .A2(n646), .ZN(n634) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n637) );
  INV_X1 U720 ( .A(n710), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n719), .ZN(n643) );
  INV_X1 U722 ( .A(KEYINPUT63), .ZN(n644) );
  XOR2_X1 U723 ( .A(G101), .B(n646), .Z(G3) );
  NAND2_X1 U724 ( .A1(n663), .A2(n648), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n647), .B(G104), .ZN(G6) );
  XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT114), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n650) );
  NAND2_X1 U728 ( .A1(n648), .A2(n665), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n652), .B(n651), .ZN(G9) );
  XOR2_X1 U731 ( .A(n653), .B(G110), .Z(G12) );
  NOR2_X1 U732 ( .A1(n660), .A2(n654), .ZN(n658) );
  XOR2_X1 U733 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n656) );
  XNOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n658), .B(n657), .ZN(G30) );
  XNOR2_X1 U737 ( .A(G143), .B(n659), .ZN(G45) );
  OR2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n662), .B(G146), .ZN(G48) );
  NAND2_X1 U740 ( .A1(n663), .A2(n666), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n664), .B(G113), .ZN(G15) );
  XOR2_X1 U742 ( .A(G116), .B(KEYINPUT117), .Z(n668) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n668), .B(n667), .ZN(G18) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT37), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  XNOR2_X1 U747 ( .A(G125), .B(n671), .ZN(G27) );
  XOR2_X1 U748 ( .A(G134), .B(n672), .Z(G36) );
  XNOR2_X1 U749 ( .A(G140), .B(n673), .ZN(G42) );
  OR2_X1 U750 ( .A1(n435), .A2(n690), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n674), .B(KEYINPUT120), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n718), .A2(n711), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(n706) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(KEYINPUT49), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n681), .Z(n682) );
  NAND2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U758 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U761 ( .A1(n690), .A2(n689), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n435), .A2(n698), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U769 ( .A(KEYINPUT119), .B(n704), .Z(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n750), .A2(n707), .ZN(n708) );
  XOR2_X1 U772 ( .A(KEYINPUT53), .B(n708), .Z(G75) );
  INV_X1 U773 ( .A(G210), .ZN(n709) );
  AND2_X1 U774 ( .A1(n711), .A2(n370), .ZN(n712) );
  NAND2_X1 U775 ( .A1(n712), .A2(n718), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n728), .A2(n716), .ZN(n717) );
  XNOR2_X1 U777 ( .A(KEYINPUT56), .B(n717), .ZN(G51) );
  NAND2_X1 U778 ( .A1(n725), .A2(G469), .ZN(n720) );
  NOR2_X1 U779 ( .A1(n728), .A2(n721), .ZN(G54) );
  XNOR2_X1 U780 ( .A(n727), .B(n726), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(KEYINPUT122), .ZN(G66) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n732) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n733), .A2(G898), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n734), .A2(n750), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n746) );
  XOR2_X1 U788 ( .A(n737), .B(KEYINPUT125), .Z(n738) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U790 ( .A(G101), .B(n740), .Z(n741) );
  NOR2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U792 ( .A(KEYINPUT124), .B(n743), .Z(n744) );
  XOR2_X1 U793 ( .A(KEYINPUT126), .B(n744), .Z(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(G69) );
  XNOR2_X1 U795 ( .A(n748), .B(n747), .ZN(n752) );
  XNOR2_X1 U796 ( .A(n749), .B(n752), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U798 ( .A(G227), .B(n752), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U802 ( .A(n757), .B(G122), .Z(G24) );
  XOR2_X1 U803 ( .A(n758), .B(G119), .Z(G21) );
  XOR2_X1 U804 ( .A(G137), .B(n759), .Z(n760) );
  XNOR2_X1 U805 ( .A(KEYINPUT127), .B(n760), .ZN(G39) );
  XNOR2_X1 U806 ( .A(n761), .B(G131), .ZN(G33) );
endmodule

