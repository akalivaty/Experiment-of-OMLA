//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n208), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n207), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n206), .B(new_n215), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n222), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT13), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  AND2_X1   g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OR2_X1    g0053(.A1(G41), .A2(G45), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n222), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT70), .B(G1698), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G226), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n257), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n250), .A2(new_n251), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT68), .A2(G1), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT68), .A2(G1), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(new_n254), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n253), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT68), .A2(G1), .ZN(new_n278));
  AND4_X1   g0078(.A1(new_n271), .A2(new_n254), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(G238), .B(new_n268), .C1(new_n275), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n248), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n258), .A2(KEYINPUT70), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G226), .ZN(new_n285));
  INV_X1    g0085(.A(new_n259), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n266), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n257), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n269), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND4_X1   g0089(.A1(new_n248), .A2(new_n280), .A3(new_n289), .A4(new_n255), .ZN(new_n290));
  OAI21_X1  g0090(.A(G169), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n280), .A2(new_n289), .A3(new_n255), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n270), .A2(new_n248), .A3(new_n280), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(G179), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT14), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(G169), .C1(new_n281), .C2(new_n290), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n277), .A2(G13), .A3(G20), .A4(new_n278), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n208), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n272), .A2(new_n273), .A3(new_n213), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n212), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n303), .B1(new_n208), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n213), .A2(new_n262), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n310), .A2(new_n217), .B1(new_n213), .B2(G68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n213), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n306), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT11), .Z(new_n316));
  NOR2_X1   g0116(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n299), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT3), .B(G33), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n260), .A3(G222), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G223), .B1(G77), .B2(new_n266), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n268), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n268), .B1(new_n275), .B2(new_n279), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n255), .B1(new_n328), .B2(new_n218), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n330), .B2(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G50), .A2(G58), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n213), .B1(new_n336), .B2(new_n208), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n338), .A2(new_n312), .B1(new_n339), .B2(new_n310), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(KEYINPUT72), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(KEYINPUT72), .B2(new_n340), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n306), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n300), .A2(G50), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G50), .B2(new_n307), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT9), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n346), .B(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT10), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n346), .B(KEYINPUT9), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT10), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n332), .A3(new_n334), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n294), .A2(new_n295), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n317), .C1(new_n356), .C2(new_n354), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n330), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n346), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(KEYINPUT73), .A2(G107), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT73), .A2(G107), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n266), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n263), .A2(new_n265), .A3(new_n282), .A4(new_n284), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n367), .B2(new_n222), .C1(new_n219), .C2(new_n324), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n256), .B1(new_n368), .B2(new_n269), .ZN(new_n369));
  OAI211_X1 g0169(.A(G244), .B(new_n268), .C1(new_n275), .C2(new_n279), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G200), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n301), .A2(new_n313), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n308), .B2(new_n313), .ZN(new_n375));
  INV_X1    g0175(.A(new_n338), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G20), .A2(G33), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(G20), .B2(G77), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  OR3_X1    g0180(.A1(new_n379), .A2(new_n380), .A3(new_n312), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n379), .B2(new_n312), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n375), .B1(new_n306), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(new_n373), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n371), .B2(new_n358), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n369), .A2(new_n360), .A3(new_n370), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n362), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AND4_X1   g0189(.A1(new_n319), .A2(new_n353), .A3(new_n357), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n300), .A2(new_n338), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n307), .B2(new_n338), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT81), .ZN(new_n393));
  INV_X1    g0193(.A(new_n306), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n320), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT76), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n395), .C1(new_n320), .C2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(G68), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n213), .B1(new_n209), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n377), .A2(G159), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n403), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G58), .A2(G68), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT77), .A3(new_n405), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n401), .A2(KEYINPUT78), .A3(new_n412), .A4(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n394), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT79), .B1(new_n264), .B2(G33), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(new_n262), .A3(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(new_n265), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n395), .A2(G20), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n208), .B1(new_n424), .B2(new_n396), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT80), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n393), .B1(new_n417), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n260), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n431));
  INV_X1    g0231(.A(G87), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n431), .A2(new_n266), .B1(new_n262), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n269), .ZN(new_n434));
  OAI211_X1 g0234(.A(G232), .B(new_n268), .C1(new_n275), .C2(new_n279), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n255), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n360), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(G169), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT18), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n407), .A2(new_n411), .ZN(new_n440));
  AOI21_X1  g0240(.A(G20), .B1(new_n263), .B2(new_n265), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n399), .B1(new_n441), .B2(KEYINPUT7), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n208), .B1(new_n442), .B2(new_n396), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n400), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT78), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n445));
  INV_X1    g0245(.A(new_n416), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n429), .B(new_n306), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n393), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n438), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G200), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n436), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G190), .B2(new_n436), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n447), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n390), .A2(new_n454), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n263), .A2(new_n265), .A3(new_n213), .A4(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT91), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT91), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n320), .A2(new_n467), .A3(new_n213), .A4(G87), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(G20), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n312), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n363), .A2(G20), .A3(new_n364), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(KEYINPUT23), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT22), .B1(new_n466), .B2(new_n468), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT24), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n466), .A2(new_n468), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n469), .A4(new_n476), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n306), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT92), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n274), .A2(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n394), .A3(new_n300), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n471), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT25), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n300), .B2(G107), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n490), .A2(G107), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n487), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n394), .B1(new_n479), .B2(new_n484), .ZN(new_n496));
  INV_X1    g0296(.A(new_n494), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT92), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n277), .A2(G45), .A3(new_n278), .ZN(new_n499));
  AND2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G264), .B(new_n268), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT5), .B(G41), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n252), .A2(new_n274), .A3(new_n504), .A4(G45), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G294), .ZN(new_n508));
  INV_X1    g0308(.A(G250), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n367), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n269), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n360), .B2(new_n512), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n495), .A2(new_n498), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT93), .B1(new_n512), .B2(G190), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n455), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT93), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n506), .A2(new_n511), .A3(new_n518), .A4(new_n356), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n486), .A3(new_n494), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n367), .C2(new_n219), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n320), .A2(new_n260), .A3(G238), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n523), .A4(new_n524), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n269), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n499), .A2(new_n509), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n274), .A2(G45), .A3(new_n249), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n268), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n489), .A2(new_n379), .ZN(new_n535));
  XOR2_X1   g0335(.A(KEYINPUT73), .B(G107), .Z(new_n536));
  NOR2_X1   g0336(.A1(G87), .A2(G97), .ZN(new_n537));
  NAND3_X1  g0337(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n537), .B1(new_n213), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n263), .A2(new_n265), .A3(new_n213), .A4(G68), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n312), .B2(new_n223), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n306), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n301), .A2(new_n379), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n534), .A2(new_n358), .B1(new_n535), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n530), .A2(new_n360), .A3(new_n533), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n490), .A2(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n545), .A3(new_n544), .ZN(new_n550));
  INV_X1    g0350(.A(new_n533), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n268), .B1(new_n525), .B2(KEYINPUT85), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n529), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n534), .A2(G200), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n547), .A2(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n263), .A2(new_n265), .A3(G250), .A4(G1698), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n320), .A2(new_n260), .A3(G244), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n320), .A2(new_n260), .A3(KEYINPUT4), .A4(G244), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n269), .ZN(new_n567));
  OAI211_X1 g0367(.A(G257), .B(new_n268), .C1(new_n499), .C2(new_n502), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n505), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n356), .A3(new_n570), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n263), .A2(new_n265), .A3(new_n282), .A4(new_n284), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT4), .A4(G244), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n268), .B1(new_n576), .B2(new_n562), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n455), .B1(new_n577), .B2(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n536), .B1(new_n424), .B2(new_n396), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n581));
  XNOR2_X1  g0381(.A(G97), .B(G107), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n584), .A2(new_n213), .B1(new_n313), .B2(new_n310), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n306), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT82), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n301), .A2(new_n587), .A3(new_n223), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT82), .B1(new_n300), .B2(G97), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n490), .A2(G97), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n586), .A2(new_n590), .A3(KEYINPUT83), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT83), .B1(new_n586), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n586), .A2(new_n590), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n358), .B1(new_n567), .B2(new_n570), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n577), .A2(new_n569), .A3(new_n360), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n556), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT86), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n567), .A2(G179), .A3(new_n570), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n577), .B2(new_n569), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n593), .A2(new_n579), .B1(new_n603), .B2(new_n595), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n556), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n262), .A2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n305), .A2(new_n212), .B1(G20), .B2(new_n473), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g0415(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT90), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(KEYINPUT20), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n614), .B(new_n620), .C1(new_n611), .C2(new_n612), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n488), .A2(G116), .A3(new_n394), .A4(new_n300), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n301), .A2(new_n473), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(G270), .B(new_n268), .C1(new_n499), .C2(new_n502), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n505), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n320), .A2(new_n260), .A3(G257), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n320), .A2(G264), .A3(G1698), .ZN(new_n630));
  XNOR2_X1  g0430(.A(KEYINPUT87), .B(G303), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n266), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT88), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n633), .A2(new_n634), .A3(new_n269), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n633), .B2(new_n269), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n628), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n625), .B1(new_n637), .B2(G200), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n356), .B2(new_n637), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n269), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT88), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n633), .A2(new_n634), .A3(new_n269), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n627), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n616), .B1(new_n613), .B2(new_n614), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n645));
  OAI21_X1  g0445(.A(G169), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT21), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT21), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n637), .A2(new_n648), .A3(new_n625), .A4(G169), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n643), .A2(new_n625), .A3(G179), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n639), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n464), .A2(new_n522), .A3(new_n607), .A4(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n362), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n349), .A2(KEYINPUT94), .A3(new_n352), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT94), .B1(new_n349), .B2(new_n352), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n388), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n318), .A2(new_n299), .B1(new_n357), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n454), .B1(new_n661), .B2(new_n462), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n655), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n464), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n514), .B1(new_n496), .B2(new_n497), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n650), .A2(new_n651), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n604), .A2(new_n666), .A3(new_n521), .A4(new_n556), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n546), .A2(new_n535), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n548), .C1(G169), .C2(new_n553), .ZN(new_n669));
  INV_X1    g0469(.A(new_n550), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n530), .A2(G190), .A3(new_n533), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n670), .B(new_n671), .C1(new_n455), .C2(new_n553), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n673), .B2(new_n598), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT83), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n595), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n586), .A2(new_n590), .A3(KEYINPUT83), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n556), .A2(new_n675), .A3(new_n603), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n667), .A2(new_n669), .A3(new_n674), .A4(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n663), .B1(new_n664), .B2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(KEYINPUT95), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n213), .A2(G13), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n274), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n625), .A2(new_n684), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n684), .B1(new_n625), .B2(new_n691), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n652), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n650), .A2(new_n651), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT96), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n639), .A3(new_n697), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n700), .B(new_n701), .C1(new_n696), .C2(new_n697), .ZN(new_n702));
  INV_X1    g0502(.A(new_n691), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n515), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n495), .A2(new_n498), .A3(new_n691), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n515), .A2(new_n705), .A3(new_n521), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n699), .A2(new_n702), .A3(G330), .A4(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n691), .B1(new_n650), .B2(new_n651), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n515), .A3(new_n521), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n665), .A2(new_n691), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(G399));
  NAND3_X1  g0513(.A1(new_n536), .A2(new_n473), .A3(new_n537), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n204), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n210), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n556), .A2(new_n594), .A3(new_n521), .A4(new_n598), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n515), .B2(new_n696), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n603), .A2(new_n679), .A3(new_n669), .A4(new_n672), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n724), .A2(KEYINPUT26), .B1(new_n548), .B2(new_n547), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n556), .A2(new_n675), .A3(new_n595), .A4(new_n603), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT29), .B(new_n703), .C1(new_n723), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n696), .A2(new_n515), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n726), .B(new_n725), .C1(new_n731), .C2(new_n722), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT98), .A3(KEYINPUT29), .A4(new_n703), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n667), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n680), .A2(new_n674), .A3(new_n669), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n703), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT97), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT97), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n681), .A2(new_n740), .A3(new_n703), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n734), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n607), .A2(new_n522), .A3(new_n653), .A4(new_n703), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n567), .A2(new_n553), .A3(new_n570), .ZN(new_n747));
  AND4_X1   g0547(.A1(G179), .A2(new_n506), .A3(new_n511), .A4(new_n626), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n641), .A2(new_n642), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n746), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n506), .A2(new_n511), .A3(G179), .A4(new_n626), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n642), .B2(new_n641), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n577), .A2(new_n569), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(KEYINPUT30), .A3(new_n754), .A4(new_n553), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n567), .A2(new_n570), .ZN(new_n756));
  AOI21_X1  g0556(.A(G179), .B1(new_n506), .B2(new_n511), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(new_n534), .A4(new_n637), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n759), .B2(new_n691), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n744), .B1(new_n745), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n743), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n743), .A2(KEYINPUT99), .A3(new_n765), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n721), .B1(new_n770), .B2(G1), .ZN(G364));
  NAND2_X1  g0571(.A1(new_n699), .A2(new_n702), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n744), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n699), .A2(new_n702), .A3(G330), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n253), .B1(new_n685), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n717), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n773), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n700), .B(new_n782), .C1(new_n696), .C2(new_n697), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n320), .A2(new_n204), .ZN(new_n784));
  INV_X1    g0584(.A(G355), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G116), .B2(new_n204), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n246), .A2(G45), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n210), .A2(G45), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(new_n716), .A3(new_n320), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n212), .B1(G20), .B2(new_n358), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n782), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n777), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n213), .A2(G190), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(G179), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(G317), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(KEYINPUT33), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(KEYINPUT33), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n213), .A2(new_n356), .A3(new_n455), .A4(G179), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G179), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n800), .B(new_n804), .C1(G329), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n213), .A2(new_n360), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n356), .A3(new_n455), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n266), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(G190), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n455), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G326), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n813), .A2(G200), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n213), .B1(new_n805), .B2(G190), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n816), .A2(G322), .B1(G294), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n795), .A2(new_n360), .A3(G200), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G283), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n808), .A2(new_n815), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n802), .A2(new_n432), .ZN(new_n824));
  OR3_X1    g0624(.A1(new_n824), .A2(KEYINPUT102), .A3(new_n266), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT102), .B1(new_n824), .B2(new_n266), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n821), .A2(G107), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT104), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n807), .A2(G159), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G50), .A2(new_n814), .B1(new_n816), .B2(G58), .ZN(new_n833));
  INV_X1    g0633(.A(new_n810), .ZN(new_n834));
  INV_X1    g0634(.A(new_n796), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G77), .A2(new_n834), .B1(new_n835), .B2(G68), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n817), .A2(new_n223), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n830), .B2(new_n831), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n833), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n823), .B1(new_n829), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n794), .B1(new_n840), .B2(new_n791), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n783), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n779), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  AND2_X1   g0644(.A1(new_n383), .A2(new_n306), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n691), .B1(new_n845), .B2(new_n375), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n385), .A2(new_n846), .B1(new_n387), .B2(new_n386), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n386), .A2(new_n387), .A3(new_n703), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT108), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT108), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n373), .A2(new_n384), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n455), .B1(new_n369), .B2(new_n370), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n388), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n855), .B2(new_n848), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n681), .A2(new_n857), .A3(new_n703), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n738), .A2(new_n741), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT108), .B1(new_n847), .B2(new_n849), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n851), .A3(new_n848), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT109), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n777), .B1(new_n865), .B2(new_n765), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n765), .B2(new_n865), .ZN(new_n867));
  INV_X1    g0667(.A(new_n791), .ZN(new_n868));
  AOI22_X1  g0668(.A1(G159), .A2(new_n834), .B1(new_n835), .B2(G150), .ZN(new_n869));
  INV_X1    g0669(.A(G137), .ZN(new_n870));
  INV_X1    g0670(.A(new_n814), .ZN(new_n871));
  INV_X1    g0671(.A(G143), .ZN(new_n872));
  INV_X1    g0672(.A(new_n816), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n869), .B1(new_n870), .B2(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT34), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n821), .A2(G68), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n807), .A2(G132), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n320), .C1(new_n802), .C2(new_n217), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(G58), .B2(new_n818), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n796), .A2(KEYINPUT105), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n796), .A2(KEYINPUT105), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(G283), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n885), .A2(new_n886), .B1(new_n473), .B2(new_n810), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n871), .A2(new_n803), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n837), .B(new_n889), .C1(G294), .C2(new_n816), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n821), .A2(G87), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n266), .B1(new_n802), .B2(new_n471), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(G311), .B2(new_n807), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n882), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n868), .B1(new_n896), .B2(KEYINPUT107), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(KEYINPUT107), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n791), .A2(new_n780), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n778), .B1(new_n313), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n898), .B(new_n900), .C1(new_n857), .C2(new_n781), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n867), .A2(new_n901), .ZN(G384));
  INV_X1    g0702(.A(new_n584), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n903), .A2(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(KEYINPUT35), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(G116), .A3(new_n214), .A4(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT36), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n211), .A2(G77), .A3(new_n403), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n217), .A2(G68), .ZN(new_n909));
  AOI211_X1 g0709(.A(G13), .B(new_n274), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n392), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n444), .A2(KEYINPUT16), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n417), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n458), .B1(new_n914), .B2(new_n689), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n438), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n449), .A2(new_n450), .ZN(new_n918));
  INV_X1    g0718(.A(new_n689), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n449), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(new_n458), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n914), .A2(new_n689), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n453), .B2(new_n462), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n858), .A2(new_n848), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n298), .A2(new_n296), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n297), .B1(new_n354), .B2(G169), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n318), .B(new_n691), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT110), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT110), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n299), .A2(new_n934), .A3(new_n318), .A4(new_n691), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n318), .A2(new_n691), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n319), .A2(new_n357), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n928), .A2(new_n940), .B1(new_n454), .B2(new_n919), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n299), .A2(new_n318), .A3(new_n703), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n458), .B1(new_n430), .B2(new_n438), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n430), .A2(new_n689), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT37), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT111), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT111), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(KEYINPUT37), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n922), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n453), .B2(new_n462), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n944), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n941), .B1(new_n943), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n734), .A2(new_n742), .A3(new_n464), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n663), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n862), .B1(new_n936), .B2(new_n938), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n760), .B1(KEYINPUT112), .B2(new_n762), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT112), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n964), .B(KEYINPUT31), .C1(new_n759), .C2(new_n691), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n745), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n967), .C1(new_n926), .C2(new_n927), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n939), .A2(new_n857), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n745), .B2(new_n966), .ZN(new_n972));
  OAI211_X1 g0772(.A(KEYINPUT40), .B(new_n972), .C1(new_n953), .C2(new_n926), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n973), .A3(new_n464), .A4(new_n967), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(G330), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n970), .A2(new_n973), .B1(new_n464), .B2(new_n967), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n961), .A2(new_n977), .B1(new_n274), .B2(new_n685), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n961), .A2(new_n977), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n911), .B1(new_n978), .B2(new_n979), .ZN(G367));
  NOR2_X1   g0780(.A1(new_n716), .A2(new_n320), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n233), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n793), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n204), .B2(new_n379), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n777), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n801), .B2(G116), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n631), .C2(new_n816), .ZN(new_n988));
  INV_X1    g0788(.A(new_n885), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(G294), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n810), .A2(new_n886), .B1(new_n820), .B2(new_n223), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n320), .B(new_n991), .C1(G317), .C2(new_n807), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n814), .A2(G311), .B1(new_n365), .B2(new_n818), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n988), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n834), .A2(G50), .B1(new_n807), .B2(G137), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n313), .B2(new_n820), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n266), .B(new_n996), .C1(G58), .C2(new_n801), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n817), .A2(new_n208), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n816), .B2(G150), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n872), .B2(new_n871), .ZN(new_n1000));
  INV_X1    g0800(.A(G159), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n997), .B1(KEYINPUT118), .B2(new_n1000), .C1(new_n1001), .C2(new_n885), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1000), .A2(KEYINPUT118), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n985), .B1(new_n1005), .B2(new_n791), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n556), .B1(new_n670), .B2(new_n703), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n547), .A2(new_n548), .A3(new_n550), .A4(new_n691), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n782), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT116), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n603), .A2(new_n679), .A3(new_n691), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n679), .A2(new_n691), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n594), .A2(new_n1014), .A3(new_n598), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT114), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n594), .A2(new_n1014), .A3(new_n598), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1013), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n710), .A2(new_n711), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1019), .A2(KEYINPUT44), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT44), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n708), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1017), .B1(new_n604), .B2(new_n1014), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1018), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1012), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n712), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1023), .A2(new_n1024), .A3(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1027), .B2(new_n712), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1019), .A2(KEYINPUT44), .A3(new_n1020), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n708), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n710), .B1(new_n707), .B2(new_n709), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n774), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n768), .A2(new_n769), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n717), .B(KEYINPUT41), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n1011), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT99), .B1(new_n743), .B2(new_n765), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n767), .B(new_n764), .C1(new_n734), .C2(new_n742), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1024), .B1(new_n1023), .B2(new_n1032), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1034), .A2(new_n1038), .A3(new_n708), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1047), .A2(new_n1048), .B1(new_n1051), .B2(new_n1042), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1045), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(KEYINPUT116), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n776), .B1(new_n1046), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT117), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1019), .A2(new_n710), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT42), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n598), .B1(new_n1019), .B2(new_n515), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n703), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT113), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(KEYINPUT43), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(KEYINPUT113), .B2(new_n1062), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1061), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1062), .A2(KEYINPUT43), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n708), .B2(new_n1019), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n708), .A2(new_n1019), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1067), .B(new_n1073), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1055), .A2(new_n1056), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1052), .A2(KEYINPUT116), .A3(new_n1053), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT116), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n775), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT117), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1010), .B1(new_n1076), .B2(new_n1081), .ZN(G387));
  INV_X1    g0882(.A(G294), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n802), .A2(new_n1083), .B1(new_n817), .B2(new_n886), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G317), .A2(new_n816), .B1(new_n834), .B2(new_n631), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT121), .B(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1085), .B1(new_n871), .B2(new_n1086), .C1(new_n885), .C2(new_n811), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT49), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n320), .B1(new_n807), .B2(G326), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n473), .C2(new_n820), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n817), .A2(new_n379), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n266), .B(new_n1094), .C1(G68), .C2(new_n834), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n802), .A2(new_n313), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n796), .A2(new_n338), .B1(new_n806), .B2(new_n339), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n821), .A2(G97), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G50), .A2(new_n816), .B1(new_n814), .B2(G159), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n868), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n715), .A2(new_n784), .B1(G107), .B2(new_n204), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n714), .B(KEYINPUT119), .Z(new_n1104));
  OR3_X1    g0904(.A1(new_n338), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT50), .B1(new_n338), .B2(G50), .ZN(new_n1106));
  AOI21_X1  g0906(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n981), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT120), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(KEYINPUT120), .B1(G45), .B2(new_n237), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1103), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n777), .B1(new_n1112), .B2(new_n793), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1102), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n782), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n707), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n770), .A2(new_n1043), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n717), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n770), .A2(new_n1043), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1116), .B1(new_n775), .B2(new_n1042), .C1(new_n1118), .C2(new_n1119), .ZN(G393));
  NAND2_X1  g0920(.A1(new_n1040), .A2(new_n776), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G150), .A2(new_n814), .B1(new_n816), .B2(G159), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT51), .Z(new_n1123));
  OAI22_X1  g0923(.A1(new_n802), .A2(new_n208), .B1(new_n810), .B2(new_n338), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n817), .A2(new_n313), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n320), .B1(new_n806), .B2(new_n872), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n989), .A2(G50), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n892), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G311), .A2(new_n816), .B1(new_n814), .B2(G317), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT52), .Z(new_n1131));
  OAI22_X1  g0931(.A1(new_n810), .A2(new_n1083), .B1(new_n806), .B2(new_n1086), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n266), .B1(new_n802), .B2(new_n886), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G116), .C2(new_n818), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n989), .A2(new_n631), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n827), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n868), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n983), .B1(new_n223), .B2(new_n204), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n243), .B2(new_n981), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1137), .A2(new_n778), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1027), .B2(new_n1115), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n717), .B1(new_n1117), .B2(new_n1051), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1040), .B1(new_n770), .B2(new_n1043), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(G390));
  NAND3_X1  g0945(.A1(new_n967), .A2(G330), .A3(new_n962), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n680), .A2(new_n674), .A3(new_n669), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n691), .B1(new_n1147), .B2(new_n667), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n849), .B1(new_n1148), .B2(new_n857), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n939), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n942), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n944), .C1(new_n953), .C2(new_n956), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n703), .B1(new_n723), .B2(new_n727), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n848), .B1(new_n1153), .B2(new_n862), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n943), .B1(new_n1154), .B2(new_n939), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n926), .B2(new_n953), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1146), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n464), .A2(G330), .A3(new_n967), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n959), .A2(new_n663), .A3(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n744), .B(new_n862), .C1(new_n745), .C2(new_n763), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1146), .B1(new_n1161), .B2(new_n939), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n929), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1154), .B1(new_n1161), .B2(new_n939), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n967), .A2(G330), .A3(new_n864), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1150), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1160), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n939), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1152), .A2(new_n1156), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1158), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT122), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n929), .A2(new_n1162), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n1160), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1160), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(KEYINPUT122), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1157), .B1(new_n1180), .B2(new_n1169), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n717), .B(new_n1171), .C1(new_n1178), .C2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n957), .A2(new_n781), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n899), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G128), .A2(new_n814), .B1(new_n816), .B2(G132), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n802), .A2(new_n339), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1187), .B2(KEYINPUT53), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n810), .A2(new_n1189), .B1(new_n820), .B2(new_n217), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n266), .B(new_n1190), .C1(G125), .C2(new_n807), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1187), .A2(KEYINPUT53), .B1(G159), .B2(new_n818), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1188), .B(new_n1193), .C1(G137), .C2(new_n989), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n871), .A2(new_n886), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1125), .B(new_n1195), .C1(G116), .C2(new_n816), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n989), .A2(new_n365), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n810), .A2(new_n223), .B1(new_n806), .B2(new_n1083), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n824), .A2(new_n320), .A3(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n878), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n777), .B1(new_n376), .B2(new_n1184), .C1(new_n1201), .C2(new_n868), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1183), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1181), .B2(new_n776), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1182), .A2(new_n1204), .ZN(G378));
  AOI21_X1  g1005(.A(new_n744), .B1(new_n968), .B2(new_n969), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n346), .A2(new_n919), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT55), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n659), .B2(new_n362), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT94), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n353), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n362), .A3(new_n656), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1210), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1208), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n659), .A2(new_n362), .A3(new_n1210), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1219), .A3(new_n1207), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1206), .A2(new_n973), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1206), .B2(new_n973), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n953), .A2(new_n956), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n923), .A2(new_n925), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT38), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n955), .B1(new_n1227), .B2(new_n954), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n943), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n940), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n954), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n453), .B2(new_n689), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1222), .A2(new_n1223), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n970), .A2(new_n973), .A3(G330), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1206), .A2(new_n973), .A3(new_n1221), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n958), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1160), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n717), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1233), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1237), .A2(new_n958), .A3(new_n1238), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n778), .B1(new_n217), .B2(new_n899), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n814), .A2(G125), .ZN(new_n1250));
  INV_X1    g1050(.A(G128), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n873), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1189), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n835), .A2(G132), .B1(new_n801), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n870), .B2(new_n810), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1252), .B(new_n1255), .C1(G150), .C2(new_n818), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G33), .A2(G41), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT123), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n820), .A2(new_n1001), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G124), .C2(new_n807), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1258), .A2(new_n1259), .A3(new_n1263), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1096), .A2(new_n998), .A3(G41), .A4(new_n320), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n471), .B2(new_n873), .C1(new_n473), .C2(new_n871), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n796), .A2(new_n223), .B1(new_n806), .B2(new_n886), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n810), .A2(new_n379), .B1(new_n820), .B2(new_n207), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(KEYINPUT58), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1261), .B(new_n217), .C1(G41), .C2(new_n320), .ZN(new_n1272));
  AND4_X1   g1072(.A1(new_n1264), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1249), .B1(new_n868), .B2(new_n1273), .C1(new_n1221), .C2(new_n781), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1246), .A2(new_n776), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1248), .A2(new_n1277), .ZN(G375));
  AOI21_X1  g1078(.A(new_n778), .B1(new_n208), .B2(new_n899), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n834), .A2(G150), .B1(new_n801), .B2(G159), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1251), .B2(new_n806), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(G132), .A2(new_n814), .B1(new_n816), .B2(G137), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n217), .B2(new_n817), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1281), .B(new_n1283), .C1(new_n989), .C2(new_n1253), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n320), .B1(new_n820), .B2(new_n207), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT126), .Z(new_n1286));
  NOR2_X1   g1086(.A1(new_n885), .A2(new_n473), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(G303), .A2(new_n807), .B1(new_n801), .B2(G97), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n266), .C1(new_n536), .C2(new_n810), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1287), .B(new_n1289), .C1(G77), .C2(new_n821), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1094), .B1(new_n814), .B2(G294), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n886), .B2(new_n873), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1284), .A2(new_n1286), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1279), .B1(new_n868), .B2(new_n1294), .C1(new_n939), .C2(new_n781), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1173), .B2(new_n775), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1173), .A2(new_n1160), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1053), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1178), .B2(new_n1299), .ZN(G381));
  OAI21_X1  g1100(.A(new_n1056), .B1(new_n1055), .B2(new_n1075), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT117), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1010), .A3(new_n1304), .ZN(new_n1305));
  OR4_X1    g1105(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1306));
  OR4_X1    g1106(.A1(G378), .A2(G375), .A3(new_n1305), .A4(new_n1306), .ZN(G407));
  AND2_X1   g1107(.A1(new_n1182), .A2(new_n1204), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n690), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G407), .B(G213), .C1(G375), .C2(new_n1309), .ZN(G409));
  OAI211_X1 g1110(.A(G378), .B(new_n1277), .C1(new_n1242), .C2(new_n1247), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1243), .A2(new_n1246), .A3(new_n1053), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1277), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G213), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(G343), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1298), .A2(KEYINPUT60), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT60), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1173), .A2(new_n1321), .A3(new_n1160), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1168), .A2(new_n718), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G384), .B1(new_n1325), .B2(new_n1297), .ZN(new_n1326));
  INV_X1    g1126(.A(G384), .ZN(new_n1327));
  AOI211_X1 g1127(.A(new_n1327), .B(new_n1296), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1317), .A2(G2897), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1326), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  AOI211_X1 g1131(.A(new_n718), .B(new_n1168), .C1(new_n1320), .C2(new_n1322), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1327), .B1(new_n1332), .B2(new_n1296), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1325), .A2(G384), .A3(new_n1297), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1331), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1317), .B1(new_n1311), .B2(new_n1314), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1338), .A2(KEYINPUT62), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT62), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1337), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(G393), .B(new_n843), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1304), .B1(new_n1303), .B2(new_n1010), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1010), .ZN(new_n1345));
  AOI211_X1 g1145(.A(new_n1345), .B(G390), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1343), .B1(new_n1344), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G387), .A2(G390), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(G393), .B(G396), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1305), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1342), .A2(new_n1351), .ZN(new_n1352));
  NOR3_X1   g1152(.A1(new_n1344), .A2(new_n1346), .A3(new_n1343), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1349), .B1(new_n1348), .B2(new_n1305), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1339), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT63), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1355), .A2(new_n1337), .A3(new_n1356), .A4(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1352), .A2(new_n1360), .ZN(G405));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1339), .A2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(G375), .A2(new_n1308), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1363), .B1(new_n1364), .B2(new_n1311), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1364), .A2(new_n1311), .A3(new_n1363), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n1355), .A3(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1367), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1351), .B1(new_n1369), .B2(new_n1365), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1368), .A2(new_n1370), .ZN(G402));
endmodule


