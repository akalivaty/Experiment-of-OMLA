

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775;

  XNOR2_X1 U369 ( .A(n485), .B(n347), .ZN(n488) );
  INV_X1 U370 ( .A(KEYINPUT16), .ZN(n347) );
  XNOR2_X1 U371 ( .A(G113), .B(G101), .ZN(n436) );
  XNOR2_X1 U372 ( .A(KEYINPUT66), .B(G131), .ZN(n452) );
  XNOR2_X2 U373 ( .A(n730), .B(n551), .ZN(n617) );
  XNOR2_X2 U374 ( .A(n550), .B(n549), .ZN(n730) );
  NAND2_X4 U375 ( .A1(n635), .A2(G953), .ZN(n666) );
  XNOR2_X2 U376 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X2 U377 ( .A(n501), .B(n351), .ZN(n508) );
  XNOR2_X2 U378 ( .A(n348), .B(G107), .ZN(n485) );
  INV_X4 U379 ( .A(G110), .ZN(n348) );
  XNOR2_X2 U380 ( .A(n583), .B(KEYINPUT38), .ZN(n725) );
  XNOR2_X2 U381 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X2 U382 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n446) );
  AND2_X2 U383 ( .A1(n381), .A2(n382), .ZN(n380) );
  NOR2_X1 U384 ( .A1(G953), .A2(G237), .ZN(n438) );
  XNOR2_X1 U385 ( .A(G113), .B(G143), .ZN(n460) );
  NAND2_X1 U386 ( .A1(G234), .A2(G237), .ZN(n430) );
  XOR2_X1 U387 ( .A(G107), .B(G122), .Z(n470) );
  NAND2_X2 U388 ( .A1(n388), .A2(n384), .ZN(n563) );
  AND2_X2 U389 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X2 U390 ( .A(G953), .ZN(n769) );
  NOR2_X1 U391 ( .A1(n742), .A2(n542), .ZN(n543) );
  OR2_X1 U392 ( .A1(n507), .A2(n534), .ZN(n542) );
  NOR2_X1 U393 ( .A1(n686), .A2(n689), .ZN(n550) );
  OR2_X1 U394 ( .A1(n477), .A2(n411), .ZN(n413) );
  AND2_X1 U395 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U396 ( .A(n397), .B(KEYINPUT35), .ZN(n774) );
  XNOR2_X1 U397 ( .A(n604), .B(KEYINPUT32), .ZN(n775) );
  XNOR2_X1 U398 ( .A(n529), .B(KEYINPUT0), .ZN(n615) );
  XNOR2_X1 U399 ( .A(n707), .B(KEYINPUT6), .ZN(n605) );
  AND2_X1 U400 ( .A1(n391), .A2(KEYINPUT106), .ZN(n377) );
  XNOR2_X1 U401 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U402 ( .A(n364), .B(n487), .ZN(n754) );
  XNOR2_X1 U403 ( .A(n363), .B(n362), .ZN(n487) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  XOR2_X1 U405 ( .A(G122), .B(G104), .Z(n486) );
  INV_X1 U406 ( .A(KEYINPUT71), .ZN(n437) );
  XNOR2_X1 U407 ( .A(G140), .B(G137), .ZN(n412) );
  NOR2_X1 U408 ( .A1(n608), .A2(n429), .ZN(n379) );
  XNOR2_X1 U409 ( .A(KEYINPUT3), .B(G116), .ZN(n362) );
  XNOR2_X1 U410 ( .A(n436), .B(G119), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U412 ( .A(n533), .B(n532), .ZN(n601) );
  XNOR2_X1 U413 ( .A(n531), .B(KEYINPUT69), .ZN(n532) );
  NAND2_X1 U414 ( .A1(n615), .A2(n374), .ZN(n533) );
  INV_X1 U415 ( .A(KEYINPUT46), .ZN(n547) );
  INV_X1 U416 ( .A(KEYINPUT44), .ZN(n373) );
  NAND2_X1 U417 ( .A1(G902), .A2(G472), .ZN(n389) );
  NAND2_X1 U418 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U419 ( .A(G472), .ZN(n387) );
  XNOR2_X1 U420 ( .A(G137), .B(KEYINPUT94), .ZN(n439) );
  XNOR2_X1 U421 ( .A(n588), .B(n587), .ZN(n354) );
  NAND2_X1 U422 ( .A1(n354), .A2(n401), .ZN(n591) );
  NOR2_X1 U423 ( .A1(n589), .A2(n402), .ZN(n401) );
  XOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n461) );
  NAND2_X1 U425 ( .A1(n489), .A2(n404), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n452), .B(G134), .ZN(n404) );
  XNOR2_X1 U427 ( .A(KEYINPUT87), .B(KEYINPUT75), .ZN(n491) );
  XOR2_X1 U428 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n492) );
  INV_X1 U429 ( .A(KEYINPUT102), .ZN(n549) );
  NOR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n444) );
  AND2_X1 U431 ( .A1(n530), .A2(n375), .ZN(n374) );
  INV_X1 U432 ( .A(n703), .ZN(n375) );
  INV_X1 U433 ( .A(KEYINPUT74), .ZN(n400) );
  NAND2_X1 U434 ( .A1(n394), .A2(n386), .ZN(n393) );
  INV_X1 U435 ( .A(G469), .ZN(n394) );
  NAND2_X1 U436 ( .A1(n670), .A2(G469), .ZN(n352) );
  XNOR2_X1 U437 ( .A(n421), .B(n420), .ZN(n647) );
  XOR2_X1 U438 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n472) );
  XNOR2_X1 U439 ( .A(KEYINPUT100), .B(KEYINPUT7), .ZN(n471) );
  XNOR2_X1 U440 ( .A(G116), .B(G134), .ZN(n469) );
  XNOR2_X1 U441 ( .A(G104), .B(G101), .ZN(n406) );
  XNOR2_X1 U442 ( .A(n488), .B(n486), .ZN(n364) );
  INV_X1 U443 ( .A(n597), .ZN(n398) );
  NOR2_X1 U444 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U445 ( .A1(n703), .A2(KEYINPUT106), .ZN(n349) );
  AND2_X1 U446 ( .A1(n354), .A2(n590), .ZN(n350) );
  NOR2_X1 U447 ( .A1(n500), .A2(n499), .ZN(n351) );
  INV_X1 U448 ( .A(G902), .ZN(n386) );
  NAND2_X1 U449 ( .A1(G902), .A2(G469), .ZN(n395) );
  INV_X1 U450 ( .A(KEYINPUT2), .ZN(n402) );
  AND2_X2 U451 ( .A1(n352), .A2(n395), .ZN(n392) );
  XNOR2_X2 U452 ( .A(n353), .B(n409), .ZN(n670) );
  XNOR2_X2 U453 ( .A(n757), .B(G146), .ZN(n353) );
  XNOR2_X1 U454 ( .A(n353), .B(n443), .ZN(n639) );
  NAND2_X2 U455 ( .A1(n356), .A2(n355), .ZN(n757) );
  OR2_X2 U456 ( .A1(n489), .A2(n404), .ZN(n356) );
  BUF_X1 U457 ( .A(n695), .Z(n357) );
  BUF_X1 U458 ( .A(n359), .Z(n707) );
  XNOR2_X1 U459 ( .A(n419), .B(n759), .ZN(n420) );
  NAND2_X1 U460 ( .A1(n380), .A2(n378), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n392), .A2(n391), .ZN(n358) );
  NAND2_X1 U462 ( .A1(n392), .A2(n391), .ZN(n506) );
  NAND2_X1 U463 ( .A1(n388), .A2(n384), .ZN(n359) );
  XNOR2_X1 U464 ( .A(n358), .B(KEYINPUT1), .ZN(n610) );
  OR2_X2 U465 ( .A1(n670), .A2(n393), .ZN(n391) );
  NOR2_X2 U466 ( .A1(n599), .A2(n703), .ZN(n608) );
  BUF_X1 U467 ( .A(n475), .Z(n479) );
  XNOR2_X1 U468 ( .A(n359), .B(KEYINPUT104), .ZN(n360) );
  XNOR2_X1 U469 ( .A(n563), .B(KEYINPUT104), .ZN(n535) );
  NAND2_X1 U470 ( .A1(n371), .A2(n373), .ZN(n369) );
  NAND2_X1 U471 ( .A1(n372), .A2(n775), .ZN(n371) );
  INV_X1 U472 ( .A(n615), .ZN(n594) );
  INV_X1 U473 ( .A(n508), .ZN(n583) );
  NAND2_X1 U474 ( .A1(n508), .A2(n724), .ZN(n562) );
  NAND2_X1 U475 ( .A1(n399), .A2(n398), .ZN(n397) );
  NOR2_X2 U476 ( .A1(n520), .A2(n516), .ZN(n686) );
  XNOR2_X1 U477 ( .A(n545), .B(KEYINPUT40), .ZN(n662) );
  XNOR2_X1 U478 ( .A(n361), .B(KEYINPUT73), .ZN(n512) );
  NAND2_X1 U479 ( .A1(n448), .A2(n449), .ZN(n361) );
  NAND2_X1 U480 ( .A1(n368), .A2(n365), .ZN(n620) );
  NAND2_X1 U481 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U482 ( .A1(n371), .A2(n373), .ZN(n366) );
  INV_X1 U483 ( .A(n598), .ZN(n367) );
  NAND2_X1 U484 ( .A1(n598), .A2(n373), .ZN(n370) );
  INV_X1 U485 ( .A(n774), .ZN(n372) );
  NAND2_X1 U486 ( .A1(n639), .A2(G472), .ZN(n390) );
  NAND2_X1 U487 ( .A1(n506), .A2(n376), .ZN(n381) );
  NOR2_X1 U488 ( .A1(n599), .A2(n349), .ZN(n376) );
  NAND2_X1 U489 ( .A1(n377), .A2(n392), .ZN(n382) );
  NAND2_X1 U490 ( .A1(n358), .A2(n608), .ZN(n383) );
  NOR2_X1 U491 ( .A1(n379), .A2(n503), .ZN(n378) );
  NOR2_X1 U492 ( .A1(n707), .A2(n383), .ZN(n614) );
  OR2_X1 U493 ( .A1(n639), .A2(n385), .ZN(n384) );
  NAND2_X1 U494 ( .A1(n535), .A2(n724), .ZN(n447) );
  XNOR2_X1 U495 ( .A(n396), .B(n400), .ZN(n449) );
  XNOR2_X1 U496 ( .A(n595), .B(n596), .ZN(n399) );
  INV_X1 U497 ( .A(n358), .ZN(n534) );
  NAND2_X1 U498 ( .A1(n610), .A2(n712), .ZN(n592) );
  INV_X1 U499 ( .A(KEYINPUT67), .ZN(n572) );
  INV_X1 U500 ( .A(KEYINPUT48), .ZN(n576) );
  INV_X1 U501 ( .A(KEYINPUT78), .ZN(n551) );
  INV_X1 U502 ( .A(KEYINPUT82), .ZN(n587) );
  INV_X1 U503 ( .A(n589), .ZN(n590) );
  INV_X1 U504 ( .A(KEYINPUT106), .ZN(n429) );
  BUF_X1 U505 ( .A(n757), .Z(n762) );
  BUF_X1 U506 ( .A(n639), .Z(n641) );
  XNOR2_X2 U507 ( .A(G143), .B(KEYINPUT77), .ZN(n403) );
  XNOR2_X2 U508 ( .A(n403), .B(G128), .ZN(n475) );
  XNOR2_X2 U509 ( .A(n475), .B(KEYINPUT4), .ZN(n489) );
  NAND2_X1 U510 ( .A1(n769), .A2(G227), .ZN(n405) );
  XNOR2_X1 U511 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U512 ( .A(n485), .B(n407), .ZN(n408) );
  XNOR2_X1 U513 ( .A(n412), .B(KEYINPUT91), .ZN(n758) );
  XNOR2_X1 U514 ( .A(n408), .B(n758), .ZN(n409) );
  NAND2_X1 U515 ( .A1(n769), .A2(G234), .ZN(n410) );
  XNOR2_X1 U516 ( .A(n410), .B(KEYINPUT8), .ZN(n477) );
  INV_X1 U517 ( .A(G221), .ZN(n411) );
  XNOR2_X1 U518 ( .A(n413), .B(n412), .ZN(n421) );
  XNOR2_X1 U519 ( .A(G119), .B(KEYINPUT23), .ZN(n415) );
  XNOR2_X1 U520 ( .A(KEYINPUT24), .B(KEYINPUT79), .ZN(n414) );
  XNOR2_X1 U521 ( .A(n415), .B(n414), .ZN(n418) );
  XNOR2_X1 U522 ( .A(G128), .B(G110), .ZN(n416) );
  XNOR2_X1 U523 ( .A(n416), .B(KEYINPUT92), .ZN(n417) );
  XNOR2_X1 U524 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U525 ( .A(G146), .B(G125), .ZN(n494) );
  XNOR2_X1 U526 ( .A(n494), .B(KEYINPUT10), .ZN(n759) );
  NAND2_X1 U527 ( .A1(n647), .A2(n386), .ZN(n426) );
  XOR2_X1 U528 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n423) );
  NAND2_X1 U529 ( .A1(n626), .A2(G234), .ZN(n422) );
  XNOR2_X1 U530 ( .A(n423), .B(n422), .ZN(n427) );
  NAND2_X1 U531 ( .A1(n427), .A2(G217), .ZN(n424) );
  XNOR2_X1 U532 ( .A(n424), .B(KEYINPUT25), .ZN(n425) );
  XNOR2_X2 U533 ( .A(n426), .B(n425), .ZN(n599) );
  NAND2_X1 U534 ( .A1(n427), .A2(G221), .ZN(n428) );
  XNOR2_X1 U535 ( .A(n428), .B(KEYINPUT21), .ZN(n703) );
  XNOR2_X1 U536 ( .A(n430), .B(KEYINPUT14), .ZN(n433) );
  NAND2_X1 U537 ( .A1(G952), .A2(n433), .ZN(n740) );
  NOR2_X1 U538 ( .A1(n740), .A2(G953), .ZN(n432) );
  INV_X1 U539 ( .A(KEYINPUT88), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n432), .B(n431), .ZN(n521) );
  NAND2_X1 U541 ( .A1(G902), .A2(n433), .ZN(n523) );
  NOR2_X1 U542 ( .A1(G900), .A2(n523), .ZN(n434) );
  NAND2_X1 U543 ( .A1(n434), .A2(G953), .ZN(n435) );
  AND2_X1 U544 ( .A1(n521), .A2(n435), .ZN(n503) );
  XNOR2_X1 U545 ( .A(n438), .B(n437), .ZN(n462) );
  NAND2_X1 U546 ( .A1(n462), .A2(G210), .ZN(n441) );
  XNOR2_X1 U547 ( .A(n439), .B(KEYINPUT5), .ZN(n440) );
  XNOR2_X1 U548 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U549 ( .A(n487), .B(n442), .Z(n443) );
  XNOR2_X1 U550 ( .A(n444), .B(KEYINPUT70), .ZN(n500) );
  INV_X1 U551 ( .A(G214), .ZN(n445) );
  OR2_X1 U552 ( .A1(n500), .A2(n445), .ZN(n724) );
  XNOR2_X1 U553 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U554 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n451) );
  XNOR2_X1 U555 ( .A(G140), .B(KEYINPUT97), .ZN(n450) );
  XOR2_X1 U556 ( .A(n451), .B(n450), .Z(n456) );
  INV_X1 U557 ( .A(n456), .ZN(n455) );
  XOR2_X1 U558 ( .A(n486), .B(n452), .Z(n453) );
  XNOR2_X1 U559 ( .A(n453), .B(n759), .ZN(n457) );
  INV_X1 U560 ( .A(n457), .ZN(n454) );
  NAND2_X1 U561 ( .A1(n455), .A2(n454), .ZN(n459) );
  NAND2_X1 U562 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U563 ( .A1(n459), .A2(n458), .ZN(n466) );
  XOR2_X1 U564 ( .A(n461), .B(n460), .Z(n464) );
  NAND2_X1 U565 ( .A1(G214), .A2(n462), .ZN(n463) );
  XNOR2_X2 U566 ( .A(n466), .B(n465), .ZN(n656) );
  NAND2_X1 U567 ( .A1(n656), .A2(n386), .ZN(n468) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(G475), .ZN(n467) );
  XNOR2_X2 U569 ( .A(n468), .B(n467), .ZN(n520) );
  INV_X1 U570 ( .A(n520), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n470), .B(n469), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U573 ( .A(n474), .B(n473), .Z(n481) );
  INV_X1 U574 ( .A(G217), .ZN(n476) );
  OR2_X1 U575 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n481), .B(n480), .ZN(n665) );
  NAND2_X1 U578 ( .A1(n665), .A2(n386), .ZN(n483) );
  INV_X1 U579 ( .A(G478), .ZN(n482) );
  XNOR2_X1 U580 ( .A(n483), .B(n482), .ZN(n519) );
  INV_X1 U581 ( .A(n519), .ZN(n516) );
  NAND2_X1 U582 ( .A1(n484), .A2(n516), .ZN(n597) );
  BUF_X1 U583 ( .A(n489), .Z(n490) );
  XNOR2_X1 U584 ( .A(n492), .B(n491), .ZN(n496) );
  NAND2_X1 U585 ( .A1(n769), .A2(G224), .ZN(n493) );
  XNOR2_X1 U586 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U587 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n490), .B(n497), .ZN(n498) );
  XNOR2_X1 U589 ( .A(n754), .B(n498), .ZN(n632) );
  NAND2_X1 U590 ( .A1(n632), .A2(n626), .ZN(n501) );
  INV_X1 U591 ( .A(G210), .ZN(n499) );
  NOR2_X1 U592 ( .A1(n597), .A2(n583), .ZN(n502) );
  AND2_X1 U593 ( .A1(n512), .A2(n502), .ZN(n568) );
  XOR2_X1 U594 ( .A(G143), .B(n568), .Z(G45) );
  NOR2_X1 U595 ( .A1(n703), .A2(n503), .ZN(n504) );
  AND2_X1 U596 ( .A1(n599), .A2(n504), .ZN(n561) );
  NAND2_X1 U597 ( .A1(n360), .A2(n561), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n505), .B(KEYINPUT28), .ZN(n507) );
  INV_X1 U599 ( .A(KEYINPUT19), .ZN(n509) );
  XNOR2_X1 U600 ( .A(n562), .B(n509), .ZN(n528) );
  NOR2_X2 U601 ( .A1(n542), .A2(n528), .ZN(n682) );
  NAND2_X1 U602 ( .A1(n682), .A2(n686), .ZN(n511) );
  XOR2_X1 U603 ( .A(G146), .B(KEYINPUT113), .Z(n510) );
  XNOR2_X1 U604 ( .A(n511), .B(n510), .ZN(G48) );
  NAND2_X1 U605 ( .A1(n512), .A2(n725), .ZN(n514) );
  XOR2_X1 U606 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n513) );
  XNOR2_X1 U607 ( .A(n514), .B(n513), .ZN(n544) );
  BUF_X1 U608 ( .A(n544), .Z(n515) );
  INV_X1 U609 ( .A(n515), .ZN(n518) );
  AND2_X1 U610 ( .A1(n520), .A2(n516), .ZN(n689) );
  INV_X1 U611 ( .A(n689), .ZN(n517) );
  NOR2_X1 U612 ( .A1(n518), .A2(n517), .ZN(n589) );
  XOR2_X1 U613 ( .A(G134), .B(n589), .Z(G36) );
  NAND2_X1 U614 ( .A1(n520), .A2(n519), .ZN(n728) );
  INV_X1 U615 ( .A(n728), .ZN(n530) );
  INV_X1 U616 ( .A(n521), .ZN(n525) );
  NOR2_X1 U617 ( .A1(n769), .A2(G898), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n522), .B(KEYINPUT89), .ZN(n753) );
  NOR2_X1 U619 ( .A1(n753), .A2(n523), .ZN(n524) );
  NOR2_X1 U620 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n526), .B(KEYINPUT90), .ZN(n527) );
  NOR2_X1 U622 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U623 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n531) );
  OR2_X1 U624 ( .A1(n601), .A2(n610), .ZN(n607) );
  INV_X1 U625 ( .A(n360), .ZN(n536) );
  NAND2_X1 U626 ( .A1(n536), .A2(n599), .ZN(n537) );
  NOR2_X1 U627 ( .A1(n607), .A2(n537), .ZN(n598) );
  XOR2_X1 U628 ( .A(G110), .B(KEYINPUT111), .Z(n538) );
  XOR2_X1 U629 ( .A(n598), .B(n538), .Z(G12) );
  NAND2_X1 U630 ( .A1(n725), .A2(n724), .ZN(n731) );
  NOR2_X1 U631 ( .A1(n728), .A2(n731), .ZN(n541) );
  XNOR2_X1 U632 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n539) );
  XOR2_X1 U633 ( .A(n539), .B(KEYINPUT109), .Z(n540) );
  XNOR2_X1 U634 ( .A(n541), .B(n540), .ZN(n742) );
  XOR2_X1 U635 ( .A(KEYINPUT42), .B(n543), .Z(n546) );
  XNOR2_X1 U636 ( .A(n546), .B(G137), .ZN(G39) );
  NAND2_X1 U637 ( .A1(n544), .A2(n686), .ZN(n545) );
  NAND2_X1 U638 ( .A1(n662), .A2(n546), .ZN(n548) );
  XNOR2_X1 U639 ( .A(n548), .B(n547), .ZN(n575) );
  INV_X1 U640 ( .A(KEYINPUT65), .ZN(n552) );
  NOR2_X1 U641 ( .A1(n617), .A2(n552), .ZN(n554) );
  NAND2_X1 U642 ( .A1(n730), .A2(KEYINPUT47), .ZN(n553) );
  NOR2_X1 U643 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U644 ( .A1(n555), .A2(n682), .ZN(n560) );
  NOR2_X1 U645 ( .A1(n617), .A2(KEYINPUT65), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n556), .A2(n682), .ZN(n558) );
  INV_X1 U647 ( .A(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U649 ( .A1(n560), .A2(n559), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n686), .A2(n561), .ZN(n578) );
  NOR2_X1 U651 ( .A1(n578), .A2(n562), .ZN(n565) );
  INV_X1 U652 ( .A(n605), .ZN(n564) );
  NAND2_X1 U653 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U654 ( .A(KEYINPUT36), .B(n566), .Z(n567) );
  NAND2_X1 U655 ( .A1(n567), .A2(n610), .ZN(n693) );
  INV_X1 U656 ( .A(n568), .ZN(n569) );
  AND2_X1 U657 ( .A1(n693), .A2(n569), .ZN(n570) );
  AND2_X1 U658 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U661 ( .A(n577), .B(n576), .ZN(n586) );
  OR2_X1 U662 ( .A1(n578), .A2(n610), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n579), .A2(n605), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n580), .A2(n724), .ZN(n581) );
  XNOR2_X1 U665 ( .A(n581), .B(KEYINPUT43), .ZN(n582) );
  XNOR2_X1 U666 ( .A(n582), .B(KEYINPUT105), .ZN(n584) );
  NOR2_X1 U667 ( .A1(n584), .A2(n508), .ZN(n694) );
  INV_X1 U668 ( .A(n694), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U670 ( .A(n591), .B(KEYINPUT81), .ZN(n622) );
  XNOR2_X1 U671 ( .A(KEYINPUT68), .B(KEYINPUT34), .ZN(n596) );
  OR2_X1 U672 ( .A1(n599), .A2(n703), .ZN(n710) );
  INV_X1 U673 ( .A(n710), .ZN(n712) );
  NOR2_X1 U674 ( .A1(n592), .A2(n605), .ZN(n593) );
  XNOR2_X1 U675 ( .A(n593), .B(KEYINPUT33), .ZN(n741) );
  NOR2_X1 U676 ( .A1(n741), .A2(n594), .ZN(n595) );
  INV_X1 U677 ( .A(n610), .ZN(n714) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT103), .ZN(n702) );
  NOR2_X1 U679 ( .A1(n714), .A2(n702), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT76), .B(n605), .Z(n600) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n702), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n676) );
  AND2_X1 U684 ( .A1(n707), .A2(n608), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT95), .ZN(n719) );
  NAND2_X1 U687 ( .A1(n615), .A2(n719), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT96), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT31), .B(n613), .ZN(n690) );
  AND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n678) );
  NOR2_X1 U691 ( .A1(n690), .A2(n678), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n676), .A2(n618), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X2 U695 ( .A(n621), .B(KEYINPUT45), .ZN(n697) );
  NAND2_X1 U696 ( .A1(n622), .A2(n697), .ZN(n624) );
  INV_X1 U697 ( .A(KEYINPUT72), .ZN(n623) );
  XNOR2_X2 U698 ( .A(n624), .B(n623), .ZN(n695) );
  NAND2_X1 U699 ( .A1(n350), .A2(n697), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n625), .A2(n402), .ZN(n628) );
  INV_X1 U701 ( .A(n626), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X4 U703 ( .A1(n695), .A2(n629), .ZN(n668) );
  NAND2_X1 U704 ( .A1(n668), .A2(G210), .ZN(n634) );
  XNOR2_X1 U705 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n630) );
  XOR2_X1 U706 ( .A(n630), .B(KEYINPUT55), .Z(n631) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n636) );
  INV_X1 U708 ( .A(G952), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n666), .ZN(n638) );
  INV_X1 U710 ( .A(KEYINPUT56), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G51) );
  NAND2_X1 U712 ( .A1(n668), .A2(G472), .ZN(n643) );
  XOR2_X1 U713 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n640) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n644), .A2(n666), .ZN(n646) );
  XNOR2_X1 U716 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(G57) );
  NAND2_X1 U718 ( .A1(n668), .A2(G217), .ZN(n649) );
  XOR2_X1 U719 ( .A(n647), .B(KEYINPUT121), .Z(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n650), .A2(n666), .ZN(n652) );
  INV_X1 U722 ( .A(KEYINPUT122), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G66) );
  NAND2_X1 U724 ( .A1(n668), .A2(G475), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT120), .B(KEYINPUT85), .Z(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT59), .B(KEYINPUT119), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n659), .A2(n666), .ZN(n661) );
  INV_X1 U730 ( .A(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(G60) );
  BUF_X1 U732 ( .A(n662), .Z(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(G131), .ZN(G33) );
  AND2_X1 U734 ( .A1(n668), .A2(G478), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n667) );
  INV_X1 U736 ( .A(n666), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n667), .A2(n674), .ZN(G63) );
  BUF_X1 U738 ( .A(n668), .Z(n669) );
  NAND2_X1 U739 ( .A1(n669), .A2(G469), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n671) );
  XNOR2_X1 U741 ( .A(n670), .B(n671), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(G54) );
  XOR2_X1 U744 ( .A(G101), .B(n676), .Z(G3) );
  NAND2_X1 U745 ( .A1(n678), .A2(n686), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(G104), .ZN(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n680) );
  NAND2_X1 U748 ( .A1(n678), .A2(n689), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U750 ( .A(G107), .B(n681), .ZN(G9) );
  NAND2_X1 U751 ( .A1(n682), .A2(n689), .ZN(n684) );
  XOR2_X1 U752 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n683) );
  XNOR2_X1 U753 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U754 ( .A(G128), .B(n685), .ZN(G30) );
  NAND2_X1 U755 ( .A1(n690), .A2(n686), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT114), .ZN(n688) );
  XNOR2_X1 U757 ( .A(G113), .B(n688), .ZN(G15) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U759 ( .A(n691), .B(G116), .ZN(G18) );
  XOR2_X1 U760 ( .A(G125), .B(KEYINPUT37), .Z(n692) );
  XNOR2_X1 U761 ( .A(n693), .B(n692), .ZN(G27) );
  XOR2_X1 U762 ( .A(G140), .B(n694), .Z(G42) );
  INV_X1 U763 ( .A(n357), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n350), .A2(KEYINPUT2), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n696), .B(KEYINPUT80), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n697), .A2(KEYINPUT2), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n746) );
  INV_X1 U769 ( .A(n702), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT115), .ZN(n706) );
  XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n706), .ZN(n709) );
  INV_X1 U773 ( .A(n707), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n718) );
  NAND2_X1 U775 ( .A1(n714), .A2(n710), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n711), .A2(KEYINPUT50), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n712), .A2(KEYINPUT50), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U782 ( .A(n721), .B(KEYINPUT116), .Z(n722) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n722), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n742), .A2(n723), .ZN(n737) );
  NOR2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U786 ( .A(KEYINPUT117), .B(n726), .Z(n727) );
  NOR2_X1 U787 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n729), .B(KEYINPUT118), .ZN(n734) );
  INV_X1 U789 ( .A(n730), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n735), .A2(n741), .ZN(n736) );
  NOR2_X1 U793 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n738), .B(KEYINPUT52), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n740), .A2(n739), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n747), .A2(G953), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n748), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U801 ( .A1(n697), .A2(n769), .ZN(n752) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n749) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n749), .ZN(n750) );
  NAND2_X1 U804 ( .A1(n750), .A2(G898), .ZN(n751) );
  NAND2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U807 ( .A(n756), .B(n755), .Z(G69) );
  XOR2_X1 U808 ( .A(KEYINPUT123), .B(n758), .Z(n760) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U810 ( .A(n762), .B(n761), .ZN(n765) );
  XNOR2_X1 U811 ( .A(n350), .B(n765), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n763), .A2(n769), .ZN(n764) );
  XOR2_X1 U813 ( .A(KEYINPUT124), .B(n764), .Z(n772) );
  XNOR2_X1 U814 ( .A(n765), .B(G227), .ZN(n766) );
  XNOR2_X1 U815 ( .A(n766), .B(KEYINPUT125), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n767), .A2(G900), .ZN(n768) );
  XOR2_X1 U817 ( .A(KEYINPUT126), .B(n768), .Z(n770) );
  NOR2_X1 U818 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U819 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U820 ( .A(KEYINPUT127), .B(n773), .ZN(G72) );
  XOR2_X1 U821 ( .A(G122), .B(n774), .Z(G24) );
  XNOR2_X1 U822 ( .A(G119), .B(n775), .ZN(G21) );
endmodule

