//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n522, new_n523, new_n524, new_n525, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT65), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G137), .A3(new_n461), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT66), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n470), .A2(new_n473), .A3(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n466), .A2(new_n461), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n467), .A2(G138), .A3(new_n461), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n474), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n487), .B2(new_n461), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n474), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n462), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n486), .A2(new_n488), .B1(new_n461), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  OR3_X1    g073(.A1(new_n497), .A2(KEYINPUT68), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT68), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n493), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G88), .B1(G50), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  AND2_X1   g088(.A1(new_n494), .A2(new_n496), .ZN(new_n514));
  AND2_X1   g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(G89), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT69), .ZN(G168));
  AOI22_X1  g096(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(new_n506), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n509), .A2(G90), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(G52), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(G301));
  INV_X1    g101(.A(G301), .ZN(G171));
  NAND2_X1  g102(.A1(G68), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G56), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n497), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT70), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n509), .A2(G81), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT71), .B(G43), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n510), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(new_n545), .A3(G53), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n510), .B2(G53), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n507), .A2(new_n508), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n514), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n550), .A2(new_n506), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G299));
  INV_X1    g131(.A(G168), .ZN(G286));
  NAND2_X1  g132(.A1(new_n509), .A2(G87), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n510), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  NAND3_X1  g136(.A1(new_n494), .A2(new_n496), .A3(G61), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT72), .A4(G61), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n510), .A2(G48), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n552), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n567), .A2(KEYINPUT73), .A3(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n509), .A2(G85), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n510), .A2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n506), .C2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n509), .A2(G92), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(KEYINPUT10), .B1(G54), .B2(new_n510), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n582), .B(KEYINPUT74), .Z(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n514), .A2(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT75), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n584), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n581), .B1(new_n592), .B2(G868), .ZN(G284));
  XNOR2_X1  g168(.A(G284), .B(KEYINPUT76), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G168), .B2(new_n595), .ZN(G297));
  XOR2_X1   g172(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n537), .A2(new_n595), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n584), .A2(new_n587), .A3(new_n591), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n603), .B2(new_n595), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g181(.A(KEYINPUT65), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n466), .B(new_n607), .ZN(new_n608));
  NOR3_X1   g183(.A1(new_n608), .A2(new_n462), .A3(G2105), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  AND2_X1   g187(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n613));
  NOR2_X1   g188(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n478), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n480), .A2(G135), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  OAI211_X1 g196(.A(new_n615), .B(new_n621), .C1(new_n613), .C2(new_n612), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2443), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n633), .B(new_n635), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT83), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT17), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  OAI22_X1  g223(.A1(new_n642), .A2(new_n646), .B1(new_n443), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n650), .B(new_n651), .Z(G227));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n658), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(KEYINPUT20), .A3(new_n655), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OAI221_X1 g238(.A(new_n660), .B1(KEYINPUT20), .B2(new_n661), .C1(new_n663), .C2(new_n658), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(G23), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G288), .B2(G16), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G1976), .ZN(new_n681));
  INV_X1    g256(.A(G1976), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n674), .A2(G22), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G303), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT90), .B(G1971), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  AND2_X1   g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n690));
  NAND2_X1  g265(.A1(G305), .A2(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n674), .A2(G6), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  AOI211_X1 g269(.A(KEYINPUT89), .B(new_n694), .C1(G305), .C2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT32), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n567), .A2(KEYINPUT73), .A3(G651), .ZN(new_n697));
  AOI21_X1  g272(.A(KEYINPUT73), .B1(new_n567), .B2(G651), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n697), .A2(new_n698), .A3(new_n573), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n699), .B2(new_n674), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n691), .A2(new_n690), .A3(new_n692), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n696), .A2(new_n704), .A3(G1981), .ZN(new_n705));
  AOI21_X1  g280(.A(G1981), .B1(new_n696), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n689), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT91), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n689), .B(new_n709), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n708), .A2(KEYINPUT34), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n708), .A2(new_n713), .A3(KEYINPUT34), .A4(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n696), .A2(new_n704), .ZN(new_n717));
  INV_X1    g292(.A(G1981), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n696), .A2(new_n704), .A3(G1981), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n709), .B1(new_n721), .B2(new_n689), .ZN(new_n722));
  INV_X1    g297(.A(new_n710), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n478), .A2(G119), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT88), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n480), .A2(G131), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT87), .B(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G25), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT35), .B(G1991), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G1986), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n674), .A2(G24), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G290), .B2(G16), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n734), .A2(new_n736), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n724), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT36), .B1(new_n715), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT34), .B1(new_n708), .B2(new_n710), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n747), .A2(new_n737), .A3(new_n743), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n748), .A2(new_n749), .A3(new_n712), .A4(new_n714), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n674), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n538), .B2(new_n674), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1341), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n478), .A2(G128), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G140), .ZN(new_n756));
  NOR2_X1   g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  INV_X1    g335(.A(new_n732), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n761), .A2(KEYINPUT28), .A3(G26), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT28), .B1(new_n761), .B2(G26), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n674), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n592), .B2(new_n674), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(new_n769), .B2(G1348), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n754), .B(new_n770), .C1(G1348), .C2(new_n769), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT93), .Z(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G11), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G33), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n480), .A2(G139), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n780), .C1(new_n781), .C2(new_n461), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(new_n775), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G2072), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(G2072), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n674), .A2(G20), .ZN(new_n787));
  OAI211_X1 g362(.A(KEYINPUT23), .B(new_n787), .C1(new_n555), .C2(new_n674), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT23), .B2(new_n787), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n761), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n761), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT29), .Z(new_n794));
  INV_X1    g369(.A(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT101), .Z(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n674), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n674), .B2(G21), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G171), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G5), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT99), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n797), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n799), .A2(new_n800), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  INV_X1    g384(.A(G160), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G34), .Z(new_n811));
  OAI22_X1  g386(.A1(new_n810), .A2(new_n775), .B1(new_n732), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G2084), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n794), .A2(new_n795), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n478), .A2(G129), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n480), .A2(G141), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT26), .Z(new_n821));
  NAND4_X1  g396(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n775), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT96), .B1(G29), .B2(G32), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT27), .B(G1996), .Z(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT30), .B(G28), .Z(new_n831));
  OAI22_X1  g406(.A1(new_n620), .A2(new_n761), .B1(G29), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n803), .B2(new_n804), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n761), .A2(G27), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G164), .B2(new_n761), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT100), .B(G2078), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n827), .A2(new_n828), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n807), .A2(new_n809), .A3(new_n830), .A4(new_n839), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n772), .A2(new_n774), .A3(new_n791), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n751), .A2(new_n841), .ZN(G150));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n843));
  NAND2_X1  g418(.A1(G150), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n751), .A2(KEYINPUT102), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(G311));
  AOI22_X1  g421(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n506), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n509), .A2(G93), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n510), .A2(G55), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n592), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n537), .B(new_n851), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT39), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n854), .B1(new_n859), .B2(G860), .ZN(G145));
  XNOR2_X1  g435(.A(new_n620), .B(new_n484), .ZN(new_n861));
  XOR2_X1   g436(.A(G160), .B(new_n861), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n783), .B(KEYINPUT104), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n610), .Z(new_n864));
  XNOR2_X1  g439(.A(G164), .B(new_n759), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g441(.A1(G130), .A2(new_n478), .B1(new_n480), .B2(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n870), .B(new_n871), .C1(G118), .C2(new_n461), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n730), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n822), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n864), .A2(new_n865), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n866), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n866), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n862), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n862), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT40), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n881), .A2(new_n884), .A3(new_n888), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(G395));
  NAND2_X1  g465(.A1(new_n852), .A2(new_n595), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n592), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n602), .A2(new_n555), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT41), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n603), .B(new_n857), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT105), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(KEYINPUT105), .B2(new_n897), .ZN(new_n900));
  XNOR2_X1  g475(.A(G303), .B(G288), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G290), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n900), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n891), .B1(new_n905), .B2(new_n595), .ZN(G295));
  OAI21_X1  g481(.A(new_n891), .B1(new_n905), .B2(new_n595), .ZN(G331));
  XNOR2_X1  g482(.A(new_n857), .B(G168), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G171), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n857), .B(G286), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G301), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n894), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n894), .B(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n909), .A3(new_n911), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n903), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n885), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n903), .B1(new_n913), .B2(new_n916), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT43), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n895), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n914), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n924), .A2(new_n909), .A3(new_n911), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n903), .B1(new_n926), .B2(new_n913), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n918), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n913), .ZN(new_n931));
  INV_X1    g506(.A(new_n903), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n919), .A2(new_n933), .A3(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n918), .B2(new_n920), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n936), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G40), .ZN(new_n941));
  NOR4_X1   g516(.A1(new_n470), .A2(new_n476), .A3(new_n941), .A4(new_n473), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT107), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n759), .B(G2067), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT108), .Z(new_n946));
  OR2_X1    g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n875), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n943), .A2(G1996), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n875), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n730), .B(new_n736), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n944), .ZN(new_n955));
  INV_X1    g530(.A(new_n943), .ZN(new_n956));
  XNOR2_X1  g531(.A(G290), .B(G1986), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n486), .A2(new_n488), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n491), .A2(new_n461), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n476), .ZN(new_n964));
  INV_X1    g539(.A(G125), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n469), .B1(new_n608), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G2105), .ZN(new_n967));
  INV_X1    g542(.A(new_n473), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n967), .A3(G40), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n973));
  NOR2_X1   g548(.A1(G288), .A2(new_n682), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n682), .A3(G288), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n977), .B2(KEYINPUT52), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n976), .B(new_n979), .C1(new_n973), .C2(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT50), .B1(new_n961), .B2(new_n962), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NOR3_X1   g561(.A1(G164), .A2(new_n986), .A3(G1384), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n942), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n795), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n942), .A2(new_n991), .A3(new_n939), .ZN(new_n992));
  INV_X1    g567(.A(G1971), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n995), .B2(new_n971), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n699), .A2(new_n718), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n574), .A2(new_n568), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G1981), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT49), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n972), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(KEYINPUT112), .A3(new_n972), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n971), .B1(new_n990), .B2(new_n994), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n984), .B(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n981), .A2(new_n996), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT125), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n992), .A2(new_n800), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n961), .A2(KEYINPUT50), .A3(new_n962), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n986), .B1(G164), .B2(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n813), .A3(new_n942), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n971), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT51), .B(G8), .C1(new_n1017), .C2(G286), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT121), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n971), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(KEYINPUT51), .C1(new_n1023), .C2(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1018), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1023), .B2(KEYINPUT122), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1019), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT126), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT62), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(new_n1019), .C1(new_n1025), .C2(new_n1031), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n992), .A2(G2078), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT53), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n992), .B2(G2078), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1040), .B(new_n1042), .C1(G1961), .C2(new_n989), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1037), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1032), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1035), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n1048), .B2(KEYINPUT59), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n963), .B2(new_n969), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n992), .B2(G1996), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(new_n538), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(new_n538), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1049), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT114), .B(G1956), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n988), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n554), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT116), .B1(new_n547), .B2(new_n548), .ZN(new_n1063));
  INV_X1    g638(.A(new_n548), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n546), .ZN(new_n1066));
  OAI221_X1 g641(.A(KEYINPUT117), .B1(new_n552), .B2(new_n553), .C1(new_n550), .C2(new_n506), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n1068), .B2(KEYINPUT115), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n555), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(KEYINPUT57), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n942), .A2(new_n991), .A3(new_n939), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1060), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT57), .A3(G299), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1069), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1058), .B1(new_n1015), .B2(new_n942), .ZN(new_n1080));
  AND4_X1   g655(.A1(new_n942), .A2(new_n991), .A3(new_n939), .A4(new_n1073), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1075), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1057), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1057), .B(KEYINPUT120), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1089));
  INV_X1    g664(.A(G1348), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n988), .A2(new_n1090), .B1(new_n970), .B2(new_n766), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(KEYINPUT60), .B2(new_n592), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1082), .B1(new_n602), .B2(new_n1091), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1075), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1040), .A2(KEYINPUT124), .A3(new_n1042), .ZN(new_n1099));
  XOR2_X1   g674(.A(G301), .B(KEYINPUT54), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(new_n1043), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1019), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1011), .B1(new_n1047), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1023), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1010), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT63), .B1(new_n1108), .B2(G168), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  OR2_X1    g686(.A1(G288), .A2(G1976), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1113));
  INV_X1    g688(.A(new_n997), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n972), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n981), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1111), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1109), .A2(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n958), .B1(new_n1106), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n953), .A2(new_n736), .A3(new_n731), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n759), .A2(G2067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n944), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n943), .A2(G1986), .A3(G290), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT48), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n955), .A2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n949), .A2(new_n947), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT47), .Z(new_n1130));
  NOR3_X1   g705(.A1(new_n1123), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1120), .A2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g707(.A1(new_n934), .A2(new_n935), .ZN(new_n1134));
  INV_X1    g708(.A(G227), .ZN(new_n1135));
  NAND4_X1  g709(.A1(new_n672), .A2(G319), .A3(new_n637), .A4(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g710(.A(new_n1136), .B(KEYINPUT127), .ZN(new_n1137));
  AND3_X1   g711(.A1(new_n886), .A2(new_n1134), .A3(new_n1137), .ZN(G308));
  NAND3_X1  g712(.A1(new_n886), .A2(new_n1134), .A3(new_n1137), .ZN(G225));
endmodule


