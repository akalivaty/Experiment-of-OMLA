

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  XNOR2_X1 U320 ( .A(n370), .B(KEYINPUT25), .ZN(n371) );
  XOR2_X1 U321 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n288) );
  XOR2_X1 U322 ( .A(n443), .B(n442), .Z(n289) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n290) );
  XNOR2_X1 U324 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U325 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U326 ( .A(n372), .B(n371), .ZN(n376) );
  XNOR2_X1 U327 ( .A(n463), .B(KEYINPUT48), .ZN(n464) );
  INV_X1 U328 ( .A(KEYINPUT94), .ZN(n380) );
  XNOR2_X1 U329 ( .A(n444), .B(n289), .ZN(n445) );
  XNOR2_X1 U330 ( .A(n465), .B(n464), .ZN(n526) );
  XNOR2_X1 U331 ( .A(n381), .B(n380), .ZN(n482) );
  XNOR2_X1 U332 ( .A(n446), .B(n445), .ZN(n452) );
  NOR2_X1 U333 ( .A1(n514), .A2(n483), .ZN(n447) );
  NOR2_X1 U334 ( .A1(n529), .A2(n473), .ZN(n562) );
  XNOR2_X1 U335 ( .A(n447), .B(KEYINPUT38), .ZN(n496) );
  XNOR2_X1 U336 ( .A(n474), .B(G169GAT), .ZN(n475) );
  XNOR2_X1 U337 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n476), .B(n475), .ZN(G1348GAT) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XNOR2_X1 U340 ( .A(G183GAT), .B(G176GAT), .ZN(n291) );
  XNOR2_X1 U341 ( .A(n288), .B(n291), .ZN(n292) );
  XOR2_X1 U342 ( .A(KEYINPUT19), .B(n292), .Z(n354) );
  XOR2_X1 U343 ( .A(G92GAT), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U346 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n296) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(n298), .B(n297), .Z(n303) );
  XOR2_X1 U350 ( .A(KEYINPUT87), .B(G64GAT), .Z(n300) );
  NAND2_X1 U351 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U353 ( .A(G8GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n354), .B(n304), .ZN(n308) );
  XOR2_X1 U356 ( .A(KEYINPUT21), .B(KEYINPUT80), .Z(n306) );
  XNOR2_X1 U357 ( .A(KEYINPUT81), .B(G211GAT), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(n307), .ZN(n345) );
  XNOR2_X1 U360 ( .A(n308), .B(n345), .ZN(n517) );
  XOR2_X1 U361 ( .A(KEYINPUT27), .B(n517), .Z(n374) );
  INV_X1 U362 ( .A(n374), .ZN(n330) );
  XOR2_X1 U363 ( .A(G85GAT), .B(G148GAT), .Z(n310) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U366 ( .A(G57GAT), .B(G120GAT), .Z(n312) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G113GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U370 ( .A(KEYINPUT86), .B(KEYINPUT1), .Z(n316) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U373 ( .A(KEYINPUT84), .B(n317), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n329) );
  XOR2_X1 U375 ( .A(KEYINPUT85), .B(KEYINPUT5), .Z(n321) );
  XNOR2_X1 U376 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n327) );
  XOR2_X1 U378 ( .A(G155GAT), .B(KEYINPUT2), .Z(n323) );
  XNOR2_X1 U379 ( .A(KEYINPUT3), .B(KEYINPUT82), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n336) );
  XOR2_X1 U381 ( .A(n336), .B(G162GAT), .Z(n325) );
  XOR2_X1 U382 ( .A(KEYINPUT0), .B(G127GAT), .Z(n352) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(n352), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U385 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n515) );
  NAND2_X1 U387 ( .A1(n330), .A2(n515), .ZN(n543) );
  XOR2_X1 U388 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n332) );
  XNOR2_X1 U389 ( .A(KEYINPUT79), .B(KEYINPUT24), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U391 ( .A(n333), .B(KEYINPUT23), .Z(n335) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U393 ( .A(G50GAT), .B(n425), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U395 ( .A(G218GAT), .B(G162GAT), .Z(n402) );
  XOR2_X1 U396 ( .A(n336), .B(n402), .Z(n338) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n347) );
  XNOR2_X1 U400 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n341), .B(KEYINPUT72), .ZN(n342) );
  XOR2_X1 U402 ( .A(n342), .B(G204GAT), .Z(n344) );
  XNOR2_X1 U403 ( .A(G78GAT), .B(G106GAT), .ZN(n343) );
  XOR2_X1 U404 ( .A(n344), .B(n343), .Z(n444) );
  XNOR2_X1 U405 ( .A(n444), .B(n345), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n470) );
  XNOR2_X1 U407 ( .A(n470), .B(KEYINPUT28), .ZN(n521) );
  NOR2_X1 U408 ( .A1(n543), .A2(n521), .ZN(n527) );
  XOR2_X1 U409 ( .A(n527), .B(KEYINPUT90), .Z(n365) );
  XOR2_X1 U410 ( .A(G15GAT), .B(G113GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n417) );
  XNOR2_X1 U413 ( .A(G99GAT), .B(G71GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n350), .B(G120GAT), .ZN(n439) );
  XNOR2_X1 U415 ( .A(n417), .B(n439), .ZN(n363) );
  AND2_X1 U416 ( .A1(G227GAT), .A2(G233GAT), .ZN(n357) );
  XOR2_X1 U417 ( .A(G190GAT), .B(G134GAT), .Z(n401) );
  XOR2_X1 U418 ( .A(KEYINPUT20), .B(KEYINPUT77), .Z(n351) );
  XNOR2_X1 U419 ( .A(n401), .B(n355), .ZN(n356) );
  NAND2_X1 U420 ( .A1(n357), .A2(n356), .ZN(n361) );
  INV_X1 U421 ( .A(n356), .ZN(n359) );
  INV_X1 U422 ( .A(n357), .ZN(n358) );
  NAND2_X1 U423 ( .A1(n359), .A2(n358), .ZN(n360) );
  NAND2_X1 U424 ( .A1(n361), .A2(n360), .ZN(n362) );
  XOR2_X1 U425 ( .A(n363), .B(n362), .Z(n366) );
  INV_X1 U426 ( .A(n366), .ZN(n529) );
  XNOR2_X1 U427 ( .A(n366), .B(KEYINPUT78), .ZN(n364) );
  NOR2_X1 U428 ( .A1(n365), .A2(n364), .ZN(n379) );
  AND2_X1 U429 ( .A1(n366), .A2(n517), .ZN(n368) );
  INV_X1 U430 ( .A(KEYINPUT91), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  NOR2_X1 U432 ( .A1(n470), .A2(n369), .ZN(n372) );
  XNOR2_X1 U433 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n370) );
  NAND2_X1 U434 ( .A1(n470), .A2(n529), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT26), .ZN(n567) );
  NOR2_X1 U436 ( .A1(n567), .A2(n374), .ZN(n375) );
  NOR2_X1 U437 ( .A1(n376), .A2(n375), .ZN(n377) );
  NOR2_X1 U438 ( .A1(n515), .A2(n377), .ZN(n378) );
  NOR2_X1 U439 ( .A1(n379), .A2(n378), .ZN(n381) );
  XNOR2_X1 U440 ( .A(G64GAT), .B(G57GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n382), .B(KEYINPUT13), .ZN(n431) );
  XOR2_X1 U442 ( .A(G8GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U443 ( .A(n431), .B(n424), .Z(n384) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n386) );
  XNOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT75), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U449 ( .A(n388), .B(n387), .Z(n396) );
  XOR2_X1 U450 ( .A(G155GAT), .B(G211GAT), .Z(n390) );
  XNOR2_X1 U451 ( .A(G22GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U453 ( .A(G127GAT), .B(G71GAT), .Z(n392) );
  XNOR2_X1 U454 ( .A(G15GAT), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n396), .B(n395), .Z(n579) );
  INV_X1 U458 ( .A(n579), .ZN(n560) );
  XNOR2_X1 U459 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n397), .B(G29GAT), .ZN(n398) );
  XOR2_X1 U461 ( .A(n398), .B(KEYINPUT7), .Z(n400) );
  XNOR2_X1 U462 ( .A(G50GAT), .B(KEYINPUT68), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n429) );
  XOR2_X1 U464 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U467 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n406) );
  XNOR2_X1 U468 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U470 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U471 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n409) );
  XOR2_X1 U472 ( .A(G92GAT), .B(G85GAT), .Z(n430) );
  XNOR2_X1 U473 ( .A(n409), .B(n430), .ZN(n410) );
  XNOR2_X1 U474 ( .A(G43GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(n429), .B(n413), .Z(n563) );
  XOR2_X1 U477 ( .A(KEYINPUT36), .B(n563), .Z(n582) );
  NOR2_X1 U478 ( .A1(n560), .A2(n582), .ZN(n414) );
  NAND2_X1 U479 ( .A1(n482), .A2(n414), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n415), .B(KEYINPUT99), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n416), .B(KEYINPUT37), .ZN(n514) );
  XOR2_X1 U482 ( .A(n417), .B(KEYINPUT30), .Z(n419) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U485 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n421) );
  XNOR2_X1 U486 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n569) );
  XNOR2_X1 U492 ( .A(KEYINPUT69), .B(n569), .ZN(n530) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  AND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  NAND2_X1 U495 ( .A1(n432), .A2(n433), .ZN(n437) );
  INV_X1 U496 ( .A(n432), .ZN(n435) );
  INV_X1 U497 ( .A(n433), .ZN(n434) );
  NAND2_X1 U498 ( .A1(n435), .A2(n434), .ZN(n436) );
  NAND2_X1 U499 ( .A1(n437), .A2(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n438), .B(KEYINPUT70), .ZN(n441) );
  XOR2_X1 U501 ( .A(n439), .B(KEYINPUT33), .Z(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U503 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n443) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n442) );
  NAND2_X1 U505 ( .A1(n530), .A2(n452), .ZN(n483) );
  AND2_X1 U506 ( .A1(n496), .A2(n366), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n449) );
  INV_X1 U508 ( .A(G43GAT), .ZN(n448) );
  INV_X1 U509 ( .A(KEYINPUT41), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n500) );
  NOR2_X1 U511 ( .A1(n500), .A2(n569), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  INV_X1 U513 ( .A(n563), .ZN(n553) );
  NOR2_X1 U514 ( .A1(n455), .A2(n563), .ZN(n456) );
  AND2_X1 U515 ( .A1(n456), .A2(n579), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(n290), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n582), .A2(n579), .ZN(n458) );
  XNOR2_X1 U518 ( .A(KEYINPUT45), .B(n458), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n459), .A2(n452), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n530), .A2(n460), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT64), .B(KEYINPUT110), .Z(n463) );
  NAND2_X1 U523 ( .A1(n526), .A2(n517), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n468), .A2(n515), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT65), .ZN(n566) );
  NOR2_X1 U528 ( .A1(n470), .A2(n566), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n562), .A2(n530), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n474) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT34), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT95), .B(n478), .Z(n485) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n480) );
  NAND2_X1 U537 ( .A1(n560), .A2(n553), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n501) );
  NOR2_X1 U540 ( .A1(n483), .A2(n501), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n490), .A2(n515), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n517), .A2(n490), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U546 ( .A1(n490), .A2(n366), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NAND2_X1 U549 ( .A1(n521), .A2(n490), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT98), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U553 ( .A1(n496), .A2(n515), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n517), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n498) );
  NAND2_X1 U558 ( .A1(n496), .A2(n521), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n504) );
  INV_X1 U562 ( .A(n500), .ZN(n555) );
  NAND2_X1 U563 ( .A1(n569), .A2(n555), .ZN(n513) );
  NOR2_X1 U564 ( .A1(n513), .A2(n501), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT103), .B(n502), .Z(n509) );
  NAND2_X1 U566 ( .A1(n509), .A2(n515), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U568 ( .A(n505), .B(G57GAT), .Z(G1332GAT) );
  NAND2_X1 U569 ( .A1(n517), .A2(n509), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U572 ( .A1(n509), .A2(n366), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n521), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U584 ( .A1(n522), .A2(n366), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n527), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n538), .A2(n530), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n533) );
  NAND2_X1 U595 ( .A1(n538), .A2(n555), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT111), .Z(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n538), .A2(n560), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U603 ( .A1(n538), .A2(n563), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT114), .Z(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n567), .A2(n543), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n526), .A2(n544), .ZN(n552) );
  NOR2_X1 U609 ( .A1(n569), .A2(n552), .ZN(n545) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U611 ( .A1(n500), .A2(n552), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT115), .B(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n579), .A2(n552), .ZN(n551) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  XOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U622 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(n568), .Z(n581) );
  NOR2_X1 U633 ( .A1(n581), .A2(n569), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n581), .A2(n452), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n581), .A2(n579), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

