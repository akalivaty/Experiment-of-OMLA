

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U554 ( .A(n730), .B(n729), .ZN(n744) );
  OR2_X1 U555 ( .A1(n691), .A2(n998), .ZN(n692) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n788) );
  AND2_X1 U557 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X4 U558 ( .A(G2105), .ZN(n524) );
  OR2_X2 U559 ( .A1(n717), .A2(n716), .ZN(n718) );
  INV_X2 U560 ( .A(n728), .ZN(n706) );
  NAND2_X2 U561 ( .A1(n688), .A2(n789), .ZN(n728) );
  NAND2_X1 U562 ( .A1(n898), .A2(G137), .ZN(n526) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n524), .ZN(n554) );
  NAND2_X1 U564 ( .A1(n775), .A2(n774), .ZN(n518) );
  OR2_X1 U565 ( .A1(n816), .A2(n520), .ZN(n519) );
  AND2_X1 U566 ( .A1(n1010), .A2(n829), .ZN(n520) );
  INV_X1 U567 ( .A(KEYINPUT64), .ZN(n694) );
  INV_X1 U568 ( .A(G8), .ZN(n731) );
  NOR2_X1 U569 ( .A1(n756), .A2(n731), .ZN(n732) );
  XNOR2_X1 U570 ( .A(n741), .B(KEYINPUT31), .ZN(n758) );
  INV_X1 U571 ( .A(n1015), .ZN(n774) );
  INV_X1 U572 ( .A(KEYINPUT74), .ZN(n588) );
  XNOR2_X1 U573 ( .A(n588), .B(KEYINPUT13), .ZN(n589) );
  XNOR2_X1 U574 ( .A(n590), .B(n589), .ZN(n591) );
  INV_X1 U575 ( .A(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U576 ( .A1(G651), .A2(n658), .ZN(n653) );
  AND2_X2 U577 ( .A1(n524), .A2(G2104), .ZN(n899) );
  NAND2_X1 U578 ( .A1(G101), .A2(n899), .ZN(n521) );
  XNOR2_X1 U579 ( .A(KEYINPUT23), .B(n521), .ZN(n528) );
  NOR2_X2 U580 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U581 ( .A(n523), .B(n522), .ZN(n898) );
  NAND2_X1 U582 ( .A1(G125), .A2(n554), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n531) );
  AND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n895) );
  NAND2_X1 U586 ( .A1(G113), .A2(n895), .ZN(n529) );
  XOR2_X1 U587 ( .A(KEYINPUT67), .B(n529), .Z(n530) );
  XNOR2_X2 U588 ( .A(n532), .B(KEYINPUT66), .ZN(G160) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n658) );
  INV_X1 U590 ( .A(G651), .ZN(n536) );
  NOR2_X1 U591 ( .A1(n658), .A2(n536), .ZN(n644) );
  NAND2_X1 U592 ( .A1(G72), .A2(n644), .ZN(n535) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n533) );
  XOR2_X2 U594 ( .A(KEYINPUT65), .B(n533), .Z(n645) );
  NAND2_X1 U595 ( .A1(G85), .A2(n645), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U597 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n537), .Z(n657) );
  NAND2_X1 U599 ( .A1(G60), .A2(n657), .ZN(n539) );
  NAND2_X1 U600 ( .A1(G47), .A2(n653), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U602 ( .A1(n541), .A2(n540), .ZN(G290) );
  NAND2_X1 U603 ( .A1(n657), .A2(G64), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT68), .ZN(n548) );
  XNOR2_X1 U605 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G77), .A2(n644), .ZN(n544) );
  NAND2_X1 U607 ( .A1(G90), .A2(n645), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G52), .A2(n653), .ZN(n549) );
  XNOR2_X1 U612 ( .A(KEYINPUT69), .B(n549), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U615 ( .A1(G111), .A2(n895), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G135), .A2(n898), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n554), .A2(G123), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT18), .B(n555), .Z(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n899), .A2(G99), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n951) );
  XNOR2_X1 U623 ( .A(G2096), .B(n951), .ZN(n560) );
  OR2_X1 U624 ( .A1(G2100), .A2(n560), .ZN(G156) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G82), .ZN(G220) );
  INV_X1 U627 ( .A(G120), .ZN(G236) );
  INV_X1 U628 ( .A(G69), .ZN(G235) );
  NAND2_X1 U629 ( .A1(G114), .A2(n895), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(KEYINPUT90), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n898), .A2(G138), .ZN(n562) );
  XOR2_X1 U632 ( .A(KEYINPUT91), .B(n562), .Z(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G126), .A2(n554), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G102), .A2(n899), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U637 ( .A1(n568), .A2(n567), .ZN(G164) );
  NAND2_X1 U638 ( .A1(G89), .A2(n645), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n569), .B(KEYINPUT4), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT76), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G76), .A2(n644), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(n573), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G63), .A2(n657), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G51), .A2(n653), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT7), .B(n580), .ZN(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n844) );
  NAND2_X1 U655 ( .A1(n844), .A2(G567), .ZN(n582) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U657 ( .A1(n657), .A2(G56), .ZN(n583) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n583), .Z(n592) );
  NAND2_X1 U659 ( .A1(G68), .A2(n644), .ZN(n587) );
  XOR2_X1 U660 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n585) );
  NAND2_X1 U661 ( .A1(G81), .A2(n645), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n653), .A2(G43), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n998) );
  INV_X1 U667 ( .A(n998), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n595), .A2(G860), .ZN(G153) );
  INV_X1 U669 ( .A(G171), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G66), .A2(n657), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G92), .A2(n645), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G79), .A2(n644), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G54), .A2(n653), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U677 ( .A(KEYINPUT75), .B(n600), .Z(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT15), .B(n603), .ZN(n997) );
  INV_X1 U680 ( .A(G868), .ZN(n670) );
  NAND2_X1 U681 ( .A1(n997), .A2(n670), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U683 ( .A1(G65), .A2(n657), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G53), .A2(n653), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G78), .A2(n644), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G91), .A2(n645), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n1001) );
  XNOR2_X1 U690 ( .A(n1001), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U691 ( .A(KEYINPUT78), .B(n670), .ZN(n612) );
  NOR2_X1 U692 ( .A1(G286), .A2(n612), .ZN(n614) );
  NOR2_X1 U693 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U695 ( .A(KEYINPUT79), .B(n615), .Z(G297) );
  INV_X1 U696 ( .A(G559), .ZN(n616) );
  NOR2_X1 U697 ( .A1(G860), .A2(n616), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n617), .B(KEYINPUT80), .ZN(n618) );
  NOR2_X1 U699 ( .A1(n997), .A2(n618), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT16), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n620), .B(KEYINPUT81), .ZN(G148) );
  NOR2_X1 U702 ( .A1(G868), .A2(n998), .ZN(n621) );
  XNOR2_X1 U703 ( .A(KEYINPUT82), .B(n621), .ZN(n624) );
  INV_X1 U704 ( .A(n997), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G868), .A2(n632), .ZN(n622) );
  NOR2_X1 U706 ( .A1(G559), .A2(n622), .ZN(n623) );
  NOR2_X1 U707 ( .A1(n624), .A2(n623), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G80), .A2(n644), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G93), .A2(n645), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U711 ( .A(KEYINPUT84), .B(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G67), .A2(n657), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G55), .A2(n653), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n671) );
  NAND2_X1 U716 ( .A1(n632), .A2(G559), .ZN(n668) );
  XOR2_X1 U717 ( .A(KEYINPUT83), .B(n998), .Z(n633) );
  XNOR2_X1 U718 ( .A(n668), .B(n633), .ZN(n634) );
  NOR2_X1 U719 ( .A1(G860), .A2(n634), .ZN(n635) );
  XOR2_X1 U720 ( .A(n671), .B(n635), .Z(G145) );
  NAND2_X1 U721 ( .A1(G61), .A2(n657), .ZN(n637) );
  NAND2_X1 U722 ( .A1(G86), .A2(n645), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n644), .A2(G73), .ZN(n638) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U727 ( .A(KEYINPUT85), .B(n641), .Z(n643) );
  NAND2_X1 U728 ( .A1(n653), .A2(G48), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G75), .A2(n644), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G88), .A2(n645), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n653), .A2(G50), .ZN(n648) );
  XOR2_X1 U734 ( .A(KEYINPUT86), .B(n648), .Z(n649) );
  NOR2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n657), .A2(G62), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G303) );
  NAND2_X1 U738 ( .A1(G49), .A2(n653), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G74), .A2(G651), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n658), .A2(G87), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(G288) );
  XNOR2_X1 U744 ( .A(n998), .B(G305), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n661) );
  XNOR2_X1 U746 ( .A(G299), .B(n661), .ZN(n664) );
  XOR2_X1 U747 ( .A(n671), .B(G290), .Z(n662) );
  XNOR2_X1 U748 ( .A(n662), .B(G303), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U750 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n667), .B(n666), .ZN(n911) );
  XNOR2_X1 U752 ( .A(n668), .B(n911), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(n678) );
  XNOR2_X1 U761 ( .A(KEYINPUT88), .B(n678), .ZN(G158) );
  XOR2_X1 U762 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G235), .A2(G236), .ZN(n679) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT89), .ZN(n680) );
  NOR2_X1 U766 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G108), .A2(n681), .ZN(n849) );
  NAND2_X1 U768 ( .A1(n849), .A2(G567), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U771 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G96), .A2(n684), .ZN(n848) );
  NAND2_X1 U773 ( .A1(n848), .A2(G2106), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n851) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U776 ( .A1(n851), .A2(n687), .ZN(n847) );
  NAND2_X1 U777 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G303), .ZN(G166) );
  XOR2_X1 U779 ( .A(KEYINPUT94), .B(n788), .Z(n688) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NAND2_X1 U781 ( .A1(n706), .A2(G1996), .ZN(n690) );
  INV_X1 U782 ( .A(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U783 ( .A(n690), .B(n689), .ZN(n693) );
  AND2_X1 U784 ( .A1(n728), .A2(G1341), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n695), .B(n694), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n704), .A2(n997), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(KEYINPUT102), .ZN(n703) );
  XNOR2_X1 U788 ( .A(KEYINPUT100), .B(KEYINPUT28), .ZN(n702) );
  NAND2_X1 U789 ( .A1(G1956), .A2(n728), .ZN(n697) );
  XNOR2_X1 U790 ( .A(KEYINPUT99), .B(n697), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n706), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U792 ( .A(KEYINPUT27), .B(n698), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n714) );
  NOR2_X1 U794 ( .A1(n714), .A2(n1001), .ZN(n701) );
  XOR2_X1 U795 ( .A(n702), .B(n701), .Z(n713) );
  AND2_X1 U796 ( .A1(n703), .A2(n713), .ZN(n712) );
  NOR2_X1 U797 ( .A1(n704), .A2(n997), .ZN(n705) );
  XNOR2_X1 U798 ( .A(KEYINPUT101), .B(n705), .ZN(n710) );
  INV_X1 U799 ( .A(n706), .ZN(n742) );
  NOR2_X1 U800 ( .A1(n706), .A2(G1348), .ZN(n708) );
  NOR2_X1 U801 ( .A1(G2067), .A2(n742), .ZN(n707) );
  NOR2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n719) );
  INV_X1 U805 ( .A(n713), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n1001), .A2(n714), .ZN(n715) );
  XOR2_X1 U807 ( .A(KEYINPUT103), .B(n715), .Z(n716) );
  AND2_X2 U808 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U809 ( .A(KEYINPUT29), .B(KEYINPUT104), .Z(n720) );
  XNOR2_X1 U810 ( .A(n721), .B(n720), .ZN(n727) );
  NAND2_X1 U811 ( .A1(G1961), .A2(n742), .ZN(n724) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n722) );
  XNOR2_X1 U813 ( .A(n722), .B(KEYINPUT97), .ZN(n921) );
  NAND2_X1 U814 ( .A1(n706), .A2(n921), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n737) );
  NOR2_X1 U816 ( .A1(G301), .A2(n737), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT98), .B(n725), .Z(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n759) );
  INV_X1 U819 ( .A(KEYINPUT95), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n728), .A2(G8), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n744), .ZN(n763) );
  INV_X1 U822 ( .A(n763), .ZN(n733) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n742), .ZN(n756) );
  NAND2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U826 ( .A1(G168), .A2(n735), .ZN(n736) );
  XNOR2_X1 U827 ( .A(n736), .B(KEYINPUT105), .ZN(n740) );
  NAND2_X1 U828 ( .A1(G301), .A2(n737), .ZN(n738) );
  XNOR2_X1 U829 ( .A(KEYINPUT106), .B(n738), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n742), .ZN(n743) );
  XNOR2_X1 U832 ( .A(KEYINPUT107), .B(n743), .ZN(n747) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n744), .ZN(n745) );
  NOR2_X1 U834 ( .A1(G166), .A2(n745), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  OR2_X1 U836 ( .A1(n731), .A2(n748), .ZN(n750) );
  AND2_X1 U837 ( .A1(n758), .A2(n750), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n759), .A2(n749), .ZN(n754) );
  INV_X1 U839 ( .A(n750), .ZN(n752) );
  AND2_X1 U840 ( .A1(G286), .A2(G8), .ZN(n751) );
  OR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U843 ( .A(KEYINPUT32), .B(n755), .Z(n765) );
  NAND2_X1 U844 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U845 ( .A(n757), .B(KEYINPUT96), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X2 U849 ( .A1(n765), .A2(n764), .ZN(n783) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n766) );
  XNOR2_X1 U851 ( .A(KEYINPUT108), .B(n766), .ZN(n772) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n772), .A2(n767), .ZN(n1008) );
  XNOR2_X1 U854 ( .A(KEYINPUT109), .B(n1008), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n783), .A2(n768), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  INV_X1 U857 ( .A(n744), .ZN(n784) );
  NAND2_X1 U858 ( .A1(n1002), .A2(n784), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U860 ( .A1(KEYINPUT33), .A2(n771), .ZN(n776) );
  AND2_X1 U861 ( .A1(n772), .A2(KEYINPUT33), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n784), .ZN(n775) );
  XNOR2_X1 U863 ( .A(G1981), .B(G305), .ZN(n1015) );
  OR2_X1 U864 ( .A1(n776), .A2(n518), .ZN(n780) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT24), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n778), .A2(n784), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G166), .A2(G8), .ZN(n781) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n817) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n829) );
  XNOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NAND2_X1 U876 ( .A1(G140), .A2(n898), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G104), .A2(n899), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n792) );
  XNOR2_X1 U880 ( .A(n793), .B(n792), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G116), .A2(n895), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G128), .A2(n554), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U884 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n799), .ZN(n881) );
  NOR2_X1 U887 ( .A1(n818), .A2(n881), .ZN(n948) );
  NAND2_X1 U888 ( .A1(n829), .A2(n948), .ZN(n826) );
  NAND2_X1 U889 ( .A1(G107), .A2(n895), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G131), .A2(n898), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G119), .A2(n554), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G95), .A2(n899), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n877) );
  AND2_X1 U896 ( .A1(n877), .A2(G1991), .ZN(n814) );
  NAND2_X1 U897 ( .A1(G117), .A2(n895), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G141), .A2(n898), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n899), .A2(G105), .ZN(n808) );
  XOR2_X1 U901 ( .A(KEYINPUT38), .B(n808), .Z(n809) );
  NOR2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n554), .A2(G129), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n907) );
  AND2_X1 U905 ( .A1(G1996), .A2(n907), .ZN(n813) );
  OR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n947) );
  NAND2_X1 U907 ( .A1(n947), .A2(n829), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n826), .A2(n819), .ZN(n816) );
  XNOR2_X1 U909 ( .A(G1986), .B(KEYINPUT92), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(G290), .ZN(n1010) );
  OR2_X1 U911 ( .A1(n817), .A2(n519), .ZN(n832) );
  NAND2_X1 U912 ( .A1(n818), .A2(n881), .ZN(n957) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n907), .ZN(n945) );
  INV_X1 U914 ( .A(n819), .ZN(n822) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n877), .ZN(n954) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n954), .A2(n820), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n945), .A2(n823), .ZN(n824) );
  XNOR2_X1 U920 ( .A(KEYINPUT39), .B(n824), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT110), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n957), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U926 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U927 ( .A(n834), .B(n833), .ZN(G329) );
  XNOR2_X1 U928 ( .A(G1341), .B(G2454), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n835), .B(G2430), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(G1348), .ZN(n842) );
  XOR2_X1 U931 ( .A(G2443), .B(G2427), .Z(n838) );
  XNOR2_X1 U932 ( .A(G2438), .B(G2446), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U934 ( .A(G2451), .B(G2435), .Z(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(G14), .ZN(n915) );
  XOR2_X1 U938 ( .A(KEYINPUT112), .B(n915), .Z(G401) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U945 ( .A(G108), .ZN(G238) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT113), .ZN(G261) );
  INV_X1 U949 ( .A(G261), .ZN(G325) );
  INV_X1 U950 ( .A(n851), .ZN(G319) );
  XNOR2_X1 U951 ( .A(G1981), .B(KEYINPUT41), .ZN(n861) );
  XOR2_X1 U952 ( .A(G1976), .B(G1961), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1956), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(G1971), .B(G1986), .Z(n855) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2474), .B(KEYINPUT114), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(G229) );
  XOR2_X1 U962 ( .A(G2100), .B(G2096), .Z(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT42), .B(G2678), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT43), .B(G2090), .Z(n865) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2072), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U968 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U969 ( .A(G2078), .B(G2084), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n554), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n895), .A2(G112), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G136), .A2(n898), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G100), .A2(n899), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U979 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n879) );
  XOR2_X1 U980 ( .A(G160), .B(n877), .Z(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(KEYINPUT117), .B(n880), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n881), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(n884), .B(G162), .Z(n894) );
  NAND2_X1 U986 ( .A1(G139), .A2(n898), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G103), .A2(n899), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n895), .A2(G115), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n887), .B(KEYINPUT116), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G127), .A2(n554), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n940) );
  XNOR2_X1 U995 ( .A(G164), .B(n940), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n894), .B(n893), .ZN(n909) );
  NAND2_X1 U997 ( .A1(G118), .A2(n895), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G130), .A2(n554), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n898), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(n902), .B(KEYINPUT45), .Z(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(n951), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n907), .B(n906), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G286), .B(n997), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n913), .B(G171), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1020 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1029) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n921), .B(G27), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT122), .B(n924), .ZN(n926) );
  XOR2_X1 U1025 ( .A(G1991), .B(G25), .Z(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(G2067), .B(G26), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G2072), .B(G33), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT121), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(G28), .A2(n932), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(KEYINPUT53), .ZN(n936) );
  XOR2_X1 U1034 ( .A(G2084), .B(KEYINPUT54), .Z(n934) );
  XNOR2_X1 U1035 ( .A(G34), .B(n934), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n967) );
  NAND2_X1 U1039 ( .A1(KEYINPUT55), .A2(n967), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n939), .ZN(n973) );
  XOR2_X1 U1041 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1042 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1044 ( .A(KEYINPUT50), .B(n943), .Z(n962) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1047 ( .A(KEYINPUT51), .B(n946), .Z(n950) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(G160), .B(G2084), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(KEYINPUT118), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT52), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT120), .ZN(n965) );
  INV_X1 U1060 ( .A(KEYINPUT55), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n968), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(G29), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(G29), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1027) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G19), .B(G1341), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(G1981), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G6), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n982), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G21), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G5), .B(G1961), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G1986), .B(KEYINPUT125), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n989), .B(G24), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n995), .Z(n996) );
  NOR2_X1 U1090 ( .A1(G16), .A2(n996), .ZN(n1024) );
  XOR2_X1 U1091 ( .A(G16), .B(KEYINPUT56), .Z(n1022) );
  XNOR2_X1 U1092 ( .A(G1348), .B(n997), .ZN(n1020) );
  XOR2_X1 U1093 ( .A(n998), .B(G1341), .Z(n1000) );
  XNOR2_X1 U1094 ( .A(G171), .B(G1961), .ZN(n999) );
  NAND2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(n1001), .B(G1956), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  INV_X1 U1098 ( .A(G1971), .ZN(n1004) );
  NOR2_X1 U1099 ( .A1(G166), .A2(n1004), .ZN(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(KEYINPUT123), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(G168), .B(G1966), .Z(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1016), .Z(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(n1025), .B(KEYINPUT126), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(n1029), .B(n1028), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

