//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n214), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n253), .A2(new_n255), .B1(G150), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n203), .A2(G20), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n251), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G50), .B1(new_n214), .B2(G1), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n262), .A2(new_n263), .B1(G50), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(new_n213), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(new_n274), .B2(new_n224), .ZN(new_n275));
  MUX2_X1   g0075(.A(G222), .B(G223), .S(G1698), .Z(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n268), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G33), .A3(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(new_n267), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G274), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  INV_X1    g0086(.A(new_n284), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n277), .B(new_n285), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(G200), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n265), .A2(KEYINPUT9), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n266), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n289), .A2(G179), .ZN(new_n296));
  INV_X1    g0096(.A(new_n265), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n285), .B1(new_n288), .B2(new_n225), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT66), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G232), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n274), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT3), .B(G33), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(KEYINPUT66), .A3(G232), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT67), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n274), .A2(G107), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n271), .A2(new_n273), .A3(G238), .A4(G1698), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n269), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n313), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n307), .B2(new_n309), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n311), .ZN(new_n319));
  OAI211_X1 g0119(.A(G190), .B(new_n303), .C1(new_n316), .C2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n252), .B(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n256), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n251), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n224), .B1(new_n260), .B2(G20), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n262), .A2(new_n328), .B1(G77), .B2(new_n261), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n319), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n269), .B1(new_n318), .B2(new_n311), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n302), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n320), .B(new_n330), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n303), .B1(new_n316), .B2(new_n319), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n330), .B1(new_n339), .B2(new_n298), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n301), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n286), .A2(new_n305), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n233), .A2(G1698), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n271), .A2(new_n344), .A3(new_n273), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n315), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n281), .A2(G238), .A3(new_n287), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n285), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G226), .A2(G1698), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n233), .B2(G1698), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n308), .B1(G33), .B2(G97), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n269), .B1(new_n359), .B2(new_n350), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(new_n349), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n356), .A2(new_n363), .A3(G190), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n356), .A2(new_n363), .A3(KEYINPUT72), .A4(G190), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n361), .B2(new_n362), .ZN(new_n370));
  OAI211_X1 g0170(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n353), .C2(new_n355), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n361), .B2(new_n362), .ZN(new_n373));
  INV_X1    g0173(.A(new_n355), .ZN(new_n374));
  AND4_X1   g0174(.A1(new_n372), .A2(new_n352), .A3(new_n362), .A4(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n370), .B(new_n371), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n255), .A2(G77), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n251), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT11), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n261), .A2(G68), .B1(KEYINPUT73), .B2(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g0182(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n214), .B2(G1), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n262), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n368), .A2(new_n377), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n376), .B2(G169), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n356), .A2(new_n363), .A3(G179), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n376), .A2(G169), .A3(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n387), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n272), .B2(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n270), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(new_n273), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n286), .A2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G223), .B2(G1698), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n269), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n285), .B1(new_n288), .B2(new_n233), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n273), .A3(new_n400), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n315), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n213), .B1(KEYINPUT65), .B2(new_n268), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n284), .B1(new_n413), .B2(new_n280), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G232), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n412), .A2(G190), .A3(new_n285), .A4(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n418));
  NAND2_X1  g0218(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n308), .B2(G20), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n274), .A2(new_n421), .A3(new_n214), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n218), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G58), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n218), .ZN(new_n425));
  OAI21_X1  g0225(.A(G20), .B1(new_n425), .B2(new_n201), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n256), .A2(G159), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n410), .A2(new_n431), .A3(new_n214), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G68), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n410), .B2(new_n214), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT16), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n429), .B(new_n250), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n262), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n252), .B1(new_n260), .B2(G20), .ZN(new_n439));
  INV_X1    g0239(.A(new_n261), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(new_n439), .B1(new_n440), .B2(new_n252), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n417), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n437), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(KEYINPUT80), .A3(new_n445), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n298), .B1(new_n407), .B2(new_n408), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n412), .A2(new_n337), .A3(new_n285), .A4(new_n415), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(KEYINPUT78), .A3(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n451), .A2(KEYINPUT78), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n437), .A2(new_n441), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(KEYINPUT79), .C2(KEYINPUT18), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n455), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n448), .A2(new_n449), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n343), .A2(new_n397), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT83), .B(new_n282), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT83), .B1(new_n471), .B2(new_n282), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n283), .A2(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n281), .A2(G274), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n227), .A2(G1698), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(G257), .B2(G1698), .ZN(new_n478));
  INV_X1    g0278(.A(G303), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n410), .A2(new_n478), .B1(new_n479), .B2(new_n308), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n473), .A2(new_n476), .B1(new_n315), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n483));
  AOI21_X1  g0283(.A(G41), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n474), .A2(new_n469), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n281), .B(G270), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n260), .A2(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n282), .B1(new_n465), .B2(new_n466), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(KEYINPUT87), .A3(G270), .A4(new_n281), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n481), .A2(new_n495), .A3(G190), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n214), .C1(G33), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT20), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  AOI22_X1  g0301(.A1(KEYINPUT88), .A2(new_n500), .B1(new_n501), .B2(G20), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n502), .A3(new_n250), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n500), .A2(KEYINPUT88), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n260), .A2(G33), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n261), .A2(new_n506), .A3(new_n213), .A4(new_n249), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G116), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G116), .B2(new_n440), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n496), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n334), .B1(new_n481), .B2(new_n495), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT89), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n481), .A2(new_n495), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT89), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n511), .A4(new_n496), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n298), .B1(new_n505), .B2(new_n509), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n520), .A3(KEYINPUT21), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n510), .A2(G179), .A3(new_n495), .A4(new_n481), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n515), .B2(new_n520), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n225), .A2(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n399), .A2(new_n400), .A3(new_n527), .A4(new_n273), .ZN(new_n528));
  XOR2_X1   g0328(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G250), .A2(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(KEYINPUT4), .A2(G244), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G1698), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n308), .A2(new_n533), .B1(G33), .B2(G283), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n315), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n473), .A2(new_n476), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n493), .A2(G257), .A3(new_n281), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n256), .A2(G77), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n498), .A3(G107), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n540), .B1(new_n544), .B2(new_n214), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n226), .B1(new_n420), .B2(new_n422), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n250), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  MUX2_X1   g0347(.A(new_n261), .B(new_n507), .S(G97), .Z(new_n548));
  AOI22_X1  g0348(.A1(new_n539), .A2(new_n298), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n492), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n469), .A3(new_n467), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n538), .B1(new_n553), .B2(new_n475), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n269), .B1(new_n530), .B2(new_n534), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n550), .B1(new_n556), .B2(new_n337), .ZN(new_n557));
  NOR4_X1   g0357(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT85), .A4(G179), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G238), .A2(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n225), .B2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(new_n273), .A3(new_n399), .A4(new_n400), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n269), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n281), .A2(G250), .A3(new_n490), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n475), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n475), .A2(new_n565), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n225), .A2(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G238), .B2(G1698), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n563), .B1(new_n410), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n315), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(G190), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n214), .B1(new_n347), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n220), .A2(new_n498), .A3(new_n226), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n399), .A2(new_n400), .A3(new_n214), .A4(new_n273), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n218), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n250), .B1(new_n440), .B2(new_n323), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n507), .A2(KEYINPUT86), .A3(new_n220), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT86), .B1(new_n507), .B2(new_n220), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n567), .A2(new_n573), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n250), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n323), .A2(new_n440), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n507), .A2(new_n323), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n298), .B1(new_n564), .B2(new_n566), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n568), .A2(new_n337), .A3(new_n572), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n554), .B2(new_n555), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT84), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n547), .A2(new_n548), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n556), .A2(G190), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(G200), .C1(new_n554), .C2(new_n555), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n559), .A2(new_n594), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n220), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n401), .A2(new_n214), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n214), .A2(G87), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n274), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n214), .B2(G107), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT90), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(new_n214), .A3(G33), .A4(G116), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT90), .B1(new_n563), .B2(G20), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n605), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n605), .A2(new_n615), .A3(KEYINPUT24), .A4(new_n607), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n250), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G13), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G1), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT25), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G20), .A4(new_n226), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT25), .B1(new_n261), .B2(G107), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n507), .C2(new_n226), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT91), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(G33), .A2(G294), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n221), .A2(new_n305), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G257), .B2(new_n305), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n410), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n315), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n493), .A2(G264), .A3(new_n281), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n553), .A2(new_n475), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n491), .A2(new_n492), .B1(new_n413), .B2(new_n280), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n315), .A2(new_n634), .B1(new_n641), .B2(G264), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT92), .B1(new_n642), .B2(new_n537), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n290), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n334), .B1(new_n637), .B2(new_n638), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n630), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n251), .B1(new_n616), .B2(new_n617), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n628), .B1(new_n647), .B2(new_n619), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n642), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G169), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n637), .A2(new_n638), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G179), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT93), .B1(new_n646), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n630), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  AOI21_X1  g0458(.A(G190), .B1(new_n649), .B2(new_n650), .ZN(new_n659));
  INV_X1    g0459(.A(new_n645), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n648), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n464), .A2(new_n526), .A3(new_n602), .A4(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n300), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT18), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT95), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT95), .B1(new_n454), .B2(new_n455), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n459), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT95), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(KEYINPUT18), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n395), .A2(new_n396), .B1(new_n388), .B2(new_n342), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n444), .A2(KEYINPUT80), .A3(new_n445), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT80), .B1(new_n444), .B2(new_n445), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n674), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n665), .B1(new_n679), .B2(new_n295), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n581), .A2(new_n584), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n564), .A2(new_n566), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(G190), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n571), .A2(KEYINPUT94), .A3(new_n315), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT94), .B1(new_n571), .B2(new_n315), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n568), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G200), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n589), .A2(new_n591), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n298), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n683), .A2(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n661), .A3(new_n559), .A4(new_n601), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n654), .A2(new_n524), .A3(new_n523), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n559), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n690), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n689), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n559), .B2(new_n593), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n463), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n680), .A2(new_n701), .ZN(G369));
  NAND2_X1  g0502(.A1(new_n622), .A2(new_n214), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n511), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n523), .B2(new_n524), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n526), .B2(new_n710), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT96), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n712), .A2(new_n713), .A3(G330), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n712), .B2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n646), .A2(new_n654), .A3(KEYINPUT93), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n658), .B1(new_n657), .B2(new_n661), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n648), .B2(new_n709), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n654), .A2(new_n708), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n709), .B1(new_n523), .B2(new_n524), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n654), .A2(new_n709), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n722), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n207), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n576), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n211), .B2(new_n731), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT97), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n683), .A2(new_n687), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n697), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT26), .B1(new_n738), .B2(new_n559), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT100), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n697), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n694), .A2(new_n695), .A3(new_n594), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n693), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT29), .B1(new_n744), .B2(new_n708), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n700), .A2(new_n709), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n747));
  INV_X1    g0547(.A(G330), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n526), .A2(new_n602), .A3(new_n708), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT99), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n719), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n559), .A2(new_n594), .A3(new_n601), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(new_n525), .A3(new_n519), .A4(new_n709), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT99), .B1(new_n753), .B2(new_n663), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n473), .A2(new_n476), .B1(G257), .B2(new_n641), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n682), .A2(new_n757), .A3(new_n536), .A4(new_n642), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n481), .A2(new_n495), .A3(G179), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(KEYINPUT98), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n758), .A2(new_n759), .A3(new_n756), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n481), .A2(new_n495), .B1(new_n642), .B2(new_n537), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(new_n686), .A3(new_n337), .A4(new_n539), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n708), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT31), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n760), .A3(new_n766), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n748), .B1(new_n755), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n747), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n736), .B1(new_n775), .B2(G1), .ZN(G364));
  NOR2_X1   g0576(.A1(new_n621), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n260), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n730), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n716), .B(new_n781), .C1(G330), .C2(new_n712), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n308), .A2(new_n207), .ZN(new_n783));
  INV_X1    g0583(.A(G355), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n784), .B1(G116), .B2(new_n207), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n401), .A2(new_n729), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n283), .B2(new_n212), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n247), .A2(G45), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n213), .B1(G20), .B2(new_n298), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n780), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n214), .A2(new_n337), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G190), .A3(new_n334), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G190), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n274), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(G20), .A3(new_n337), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n801), .B(new_n805), .C1(G329), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n798), .A2(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n290), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G326), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n214), .A2(new_n334), .A3(G179), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n809), .A2(G190), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G303), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n290), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n337), .A2(new_n334), .A3(G190), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n819), .A2(G283), .B1(new_n821), .B2(G294), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n808), .A2(new_n811), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n813), .A2(new_n220), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n807), .A2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(new_n815), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(KEYINPUT32), .B2(new_n826), .C1(new_n218), .C2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G107), .A2(new_n819), .B1(new_n826), .B2(KEYINPUT32), .ZN(new_n829));
  INV_X1    g0629(.A(new_n810), .ZN(new_n830));
  INV_X1    g0630(.A(new_n821), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n202), .B2(new_n830), .C1(new_n498), .C2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n308), .B1(new_n803), .B2(new_n224), .C1(new_n424), .C2(new_n799), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n823), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n797), .B1(new_n835), .B2(new_n794), .ZN(new_n836));
  INV_X1    g0636(.A(new_n793), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n712), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n782), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  OAI21_X1  g0640(.A(new_n708), .B1(new_n326), .B2(new_n329), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n335), .A2(new_n841), .B1(new_n340), .B2(new_n338), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n341), .A2(new_n708), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n746), .B(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n774), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n780), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  INV_X1    g0650(.A(new_n844), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n791), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n813), .A2(new_n226), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n818), .A2(new_n220), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(G303), .C2(new_n810), .ZN(new_n856));
  INV_X1    g0656(.A(G294), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n799), .A2(new_n857), .B1(new_n806), .B2(new_n804), .ZN(new_n858));
  INV_X1    g0658(.A(new_n803), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n308), .B(new_n858), .C1(G116), .C2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n815), .A2(G283), .B1(G97), .B2(new_n821), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n856), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n799), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(G143), .B1(new_n859), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G150), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n827), .B2(new_n865), .C1(new_n866), .C2(new_n830), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n410), .B1(G132), .B2(new_n807), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n818), .A2(new_n218), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n424), .B2(new_n831), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G50), .B2(new_n814), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n867), .A2(new_n868), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n862), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n853), .B1(new_n877), .B2(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT102), .B2(new_n877), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n853), .A2(new_n792), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n780), .B1(G77), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT101), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n849), .A2(new_n850), .B1(new_n852), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  INV_X1    g0685(.A(new_n747), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n886), .A2(KEYINPUT104), .A3(new_n464), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT104), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n747), .B2(new_n463), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n680), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n461), .A2(new_n456), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n676), .B2(new_n677), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n250), .B1(new_n435), .B2(new_n436), .ZN(new_n893));
  INV_X1    g0693(.A(new_n418), .ZN(new_n894));
  INV_X1    g0694(.A(new_n434), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G68), .A3(new_n432), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n896), .B2(new_n430), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n441), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n706), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n454), .A2(new_n898), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n900), .A3(new_n442), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n706), .B1(new_n437), .B2(new_n441), .ZN(new_n905));
  INV_X1    g0705(.A(new_n455), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n417), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT37), .B1(new_n454), .B2(new_n455), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n904), .A2(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n912), .B(new_n909), .C1(new_n892), .C2(new_n901), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n905), .ZN(new_n916));
  INV_X1    g0716(.A(new_n446), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n674), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n907), .B1(new_n667), .B2(new_n668), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n912), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT39), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n395), .A2(new_n396), .A3(new_n709), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n915), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n911), .A2(new_n913), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n844), .B(new_n709), .C1(new_n693), .C2(new_n699), .ZN(new_n927));
  INV_X1    g0727(.A(new_n843), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n396), .B(new_n708), .C1(new_n395), .C2(new_n389), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n394), .A2(new_n393), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n396), .B1(new_n931), .B2(new_n391), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n396), .A2(new_n708), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n388), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n926), .A2(new_n936), .B1(new_n674), .B2(new_n899), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n925), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n890), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n767), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n770), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n755), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n851), .B1(new_n930), .B2(new_n934), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n940), .B1(new_n946), .B2(new_n926), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n921), .A2(new_n922), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n948), .A2(KEYINPUT40), .A3(new_n944), .A4(new_n945), .ZN(new_n949));
  AND4_X1   g0749(.A1(new_n463), .A2(new_n947), .A3(new_n944), .A4(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n947), .A2(new_n949), .B1(new_n463), .B2(new_n944), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n950), .A2(new_n748), .A3(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n939), .A2(new_n952), .B1(new_n260), .B2(new_n777), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n939), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(new_n544), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT35), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT35), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n956), .A2(G116), .A3(new_n215), .A4(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT36), .Z(new_n959));
  OR3_X1    g0759(.A1(new_n211), .A2(new_n224), .A3(new_n425), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n202), .A2(G68), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT103), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n260), .B(G13), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n954), .A2(new_n959), .A3(new_n963), .ZN(G367));
  NAND2_X1  g0764(.A1(new_n814), .A2(G116), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT46), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n831), .A2(new_n226), .B1(new_n818), .B2(new_n498), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G294), .B2(new_n815), .ZN(new_n968));
  INV_X1    g0768(.A(G283), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n799), .A2(new_n479), .B1(new_n803), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G317), .B2(new_n807), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n401), .B1(new_n810), .B2(G311), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n819), .A2(G77), .ZN(new_n974));
  INV_X1    g0774(.A(G159), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n424), .B2(new_n813), .C1(new_n975), .C2(new_n827), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n821), .A2(G68), .ZN(new_n977));
  INV_X1    g0777(.A(G143), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n830), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n308), .B1(new_n806), .B2(new_n866), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n799), .A2(new_n865), .B1(new_n803), .B2(new_n202), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n973), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n794), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n796), .B1(new_n729), .B2(new_n324), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n239), .A2(new_n786), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n781), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n681), .A2(new_n708), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n690), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n697), .B2(new_n989), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n985), .B(new_n988), .C1(new_n837), .C2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n775), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT107), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n559), .A2(new_n709), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT105), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n559), .B(new_n601), .C1(new_n597), .C2(new_n709), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n727), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT44), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n726), .A3(new_n725), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n1004));
  XOR2_X1   g0804(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n722), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1001), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n722), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1003), .B(new_n1004), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n725), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n714), .B2(new_n715), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n716), .A2(new_n725), .A3(new_n1013), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n775), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n995), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1018), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1020), .A2(new_n1006), .A3(KEYINPUT107), .A4(new_n1011), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n994), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n730), .B(KEYINPUT41), .Z(new_n1023));
  OAI21_X1  g0823(.A(new_n778), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n559), .B1(new_n1000), .B2(new_n657), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n999), .A2(new_n719), .A3(new_n724), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n709), .B1(KEYINPUT42), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT42), .B2(new_n1026), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1028), .A2(KEYINPUT43), .A3(new_n991), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n722), .A2(new_n999), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1034), .B(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n993), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(G387));
  NAND3_X1  g0839(.A1(new_n720), .A2(new_n721), .A3(new_n793), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n783), .A2(new_n732), .B1(G107), .B2(new_n207), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n321), .A2(new_n202), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI21_X1  g0845(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n732), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n787), .B1(new_n236), .B2(G45), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n780), .B1(new_n1049), .B2(new_n796), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n410), .B1(G150), .B2(new_n807), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n224), .B2(new_n813), .C1(new_n498), .C2(new_n818), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT109), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n799), .A2(new_n202), .B1(new_n803), .B2(new_n218), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n831), .A2(new_n323), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n975), .B2(new_n830), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(new_n253), .C2(new_n815), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n401), .B1(G326), .B2(new_n807), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n831), .A2(new_n969), .B1(new_n813), .B2(new_n857), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n863), .A2(G317), .B1(new_n859), .B2(G303), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n827), .B2(new_n804), .C1(new_n800), .C2(new_n830), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1060), .B1(new_n501), .B2(new_n818), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1050), .B1(new_n1070), .B2(new_n794), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1017), .A2(new_n779), .B1(new_n1040), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1018), .A2(new_n730), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1017), .A2(new_n775), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(G393));
  NAND2_X1  g0875(.A1(new_n244), .A2(new_n786), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n796), .B1(G97), .B2(new_n729), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n781), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT110), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(KEYINPUT110), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G317), .A2(new_n810), .B1(new_n863), .B2(G311), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n274), .B1(new_n806), .B2(new_n800), .C1(new_n803), .C2(new_n857), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n827), .A2(new_n479), .B1(new_n226), .B2(new_n818), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n831), .A2(new_n501), .B1(new_n813), .B2(new_n969), .ZN(new_n1085));
  OR4_X1    g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n830), .A2(new_n865), .B1(new_n975), .B2(new_n799), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n827), .A2(new_n202), .B1(new_n218), .B2(new_n813), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n831), .A2(new_n224), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1089), .A2(new_n855), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n401), .B1(new_n978), .B2(new_n806), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n321), .B2(new_n859), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1080), .B1(new_n1095), .B2(new_n794), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1079), .B(new_n1096), .C1(new_n999), .C2(new_n837), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1012), .B2(new_n778), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT111), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n731), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  INV_X1    g0903(.A(new_n924), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n929), .B2(new_n935), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n667), .A2(new_n668), .A3(new_n666), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n917), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n905), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n920), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT38), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n914), .B1(new_n1111), .B2(new_n913), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n910), .B1(new_n462), .B2(new_n900), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n912), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1105), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n774), .A2(new_n844), .A3(new_n935), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n842), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n709), .B(new_n1119), .C1(new_n743), .C2(new_n693), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n928), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n935), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n948), .A2(new_n1122), .A3(new_n924), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1116), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n936), .A2(new_n924), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n915), .B2(new_n923), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n948), .A2(new_n924), .A3(new_n1122), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n779), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n791), .B1(new_n915), .B2(new_n923), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n780), .B1(new_n253), .B2(new_n880), .ZN(new_n1133));
  INV_X1    g0933(.A(G132), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n799), .A2(new_n1134), .B1(new_n803), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n274), .B(new_n1136), .C1(G125), .C2(new_n807), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n813), .A2(new_n865), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n819), .A2(G50), .B1(new_n815), .B2(G137), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n810), .A2(G128), .B1(G159), .B2(new_n821), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n799), .A2(new_n501), .B1(new_n806), .B2(new_n857), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n308), .B(new_n1143), .C1(G97), .C2(new_n859), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n825), .A3(new_n872), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1090), .B1(G283), .B2(new_n810), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n226), .B2(new_n827), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1133), .B1(new_n1148), .B2(new_n794), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1132), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1131), .A2(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT113), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n932), .A2(new_n388), .A3(new_n933), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n933), .B1(new_n932), .B2(new_n388), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n844), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n942), .B1(new_n751), .B2(new_n754), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n748), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1127), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1121), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1156), .A2(new_n748), .A3(new_n851), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1117), .B(new_n1161), .C1(new_n935), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n935), .B1(new_n774), .B2(new_n844), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n929), .B1(new_n1165), .B2(new_n1157), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT112), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n770), .A2(new_n772), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n751), .B2(new_n754), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1169), .A2(new_n748), .A3(new_n851), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1125), .B1(new_n1170), .B2(new_n935), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT112), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n929), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1164), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n463), .A2(new_n944), .A3(G330), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n680), .B(new_n1175), .C1(new_n887), .C2(new_n889), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1160), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n929), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n750), .B1(new_n749), .B2(new_n719), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n753), .A2(new_n663), .A3(KEYINPUT99), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n773), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(G330), .A3(new_n844), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n935), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(KEYINPUT112), .B(new_n1178), .C1(new_n1184), .C2(new_n1125), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1172), .B1(new_n1171), .B2(new_n929), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1163), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1176), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1130), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1177), .A2(new_n1189), .A3(new_n730), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1151), .A2(KEYINPUT113), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1152), .A2(new_n1190), .A3(new_n1191), .ZN(G378));
  NOR2_X1   g0992(.A1(new_n265), .A2(new_n706), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n301), .B(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n791), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n780), .B1(G50), .B2(new_n880), .ZN(new_n1200));
  OR3_X1    g1000(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n1135), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT116), .B1(new_n813), .B2(new_n1135), .ZN(new_n1202));
  INV_X1    g1002(.A(G128), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1202), .C1(new_n1203), .C2(new_n799), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT117), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n810), .A2(G125), .B1(new_n859), .B2(G137), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n815), .A2(G132), .B1(G150), .B2(new_n821), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT59), .Z(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n975), .C2(new_n818), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n410), .A2(new_n282), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G77), .B2(new_n814), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT115), .Z(new_n1214));
  NOR2_X1   g1014(.A1(new_n818), .A2(new_n424), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT114), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n863), .A2(G107), .B1(G283), .B2(new_n807), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n323), .B2(new_n803), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n977), .B1(new_n827), .B2(new_n498), .C1(new_n501), .C2(new_n830), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1214), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1212), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1211), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1200), .B1(new_n1225), .B2(new_n794), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT118), .B1(new_n1199), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1199), .A2(KEYINPUT118), .A3(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT119), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n947), .A2(G330), .A3(new_n949), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1198), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n947), .A2(new_n1197), .A3(G330), .A4(new_n949), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n938), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n938), .A3(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n779), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1231), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1188), .B1(new_n1174), .B2(new_n1160), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT120), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(KEYINPUT120), .B(new_n1188), .C1(new_n1174), .C2(new_n1160), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1238), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT57), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n731), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1240), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1023), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1183), .A2(new_n791), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n780), .B1(G68), .B2(new_n880), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n501), .A2(new_n827), .B1(new_n830), .B2(new_n857), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G97), .B2(new_n814), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n799), .A2(new_n969), .B1(new_n803), .B2(new_n226), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n308), .B(new_n1261), .C1(G303), .C2(new_n807), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1260), .A2(new_n974), .A3(new_n1056), .A4(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n859), .A2(G150), .B1(new_n807), .B2(G128), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n814), .A2(G159), .B1(new_n821), .B2(G50), .ZN(new_n1265));
  AND4_X1   g1065(.A1(new_n401), .A2(new_n1216), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n827), .A2(new_n1135), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G137), .B2(new_n863), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1267), .B(new_n1269), .C1(new_n1134), .C2(new_n830), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1263), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1258), .B1(new_n1272), .B2(new_n794), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1187), .A2(new_n779), .B1(new_n1257), .B2(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1256), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(G381));
  INV_X1    g1076(.A(new_n1151), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1190), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT122), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT122), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1190), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1038), .A2(new_n1102), .A3(new_n1275), .A4(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1251), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1286), .B2(new_n1251), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G213), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1283), .A2(G343), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1251), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(G409));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1236), .A2(new_n1297), .A3(new_n1237), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1233), .A2(new_n938), .A3(new_n1234), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT126), .B1(new_n1299), .B2(new_n1235), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1300), .A3(new_n779), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1255), .B1(new_n1299), .B2(new_n1235), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1230), .B(new_n1301), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  AOI211_X1 g1105(.A(KEYINPUT125), .B(new_n1302), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1282), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1240), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1176), .B1(new_n1187), .B2(new_n1130), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(KEYINPUT120), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1244), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1249), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n730), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1238), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G378), .B(new_n1308), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1291), .A2(G343), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1253), .A2(KEYINPUT60), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1254), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1176), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1324), .A2(new_n730), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(G384), .A3(new_n1274), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1326), .B2(new_n1274), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1321), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1274), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n884), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1327), .A3(new_n1320), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1336), .B1(new_n1319), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1038), .A2(G390), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1038), .A2(G390), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(G393), .B(new_n839), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(KEYINPUT127), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1343), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1344), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1347), .B1(new_n1343), .B2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1317), .B1(new_n1307), .B2(new_n1315), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1335), .A2(new_n1339), .A3(new_n1350), .A4(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT62), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1351), .A2(new_n1354), .A3(new_n1337), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT61), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1356), .B1(new_n1351), .B2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1354), .B1(new_n1351), .B2(new_n1337), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1355), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1353), .B1(new_n1360), .B2(new_n1350), .ZN(G405));
  OAI21_X1  g1161(.A(new_n1315), .B1(new_n1251), .B2(new_n1283), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1362), .B(new_n1338), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(new_n1350), .ZN(G402));
endmodule


