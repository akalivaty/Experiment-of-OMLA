//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g027(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n466), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n477), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n476), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n477), .C1(new_n463), .C2(new_n464), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G138), .A4(new_n477), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(KEYINPUT67), .B2(G114), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT67), .A2(G114), .ZN(new_n494));
  OAI211_X1 g069(.A(G2104), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT67), .A2(G114), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(G2105), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .A3(G2104), .A4(new_n492), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n491), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G50), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(new_n508), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G543), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n525), .A2(G88), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n514), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT70), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n514), .A2(new_n524), .A3(new_n528), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G166));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n513), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G63), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n507), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n509), .B2(new_n511), .ZN(new_n539));
  NOR3_X1   g114(.A1(new_n539), .A2(new_n516), .A3(new_n508), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n537), .A2(new_n527), .B1(G51), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n512), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n539), .A2(new_n508), .A3(new_n520), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G90), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT72), .B(G52), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n512), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT73), .B(G43), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n540), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT74), .B(G81), .Z(new_n558));
  NAND2_X1  g133(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(KEYINPUT75), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n557), .B2(new_n559), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n555), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  OAI211_X1 g146(.A(G543), .B(new_n526), .C1(new_n523), .C2(new_n538), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n513), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(KEYINPUT76), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n574), .B2(new_n576), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(KEYINPUT78), .A2(G65), .ZN(new_n582));
  NAND2_X1  g157(.A1(KEYINPUT78), .A2(G65), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n527), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n507), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n513), .A2(new_n587), .A3(new_n527), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n526), .B(new_n527), .C1(new_n523), .C2(new_n538), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n586), .B1(new_n591), .B2(G91), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n581), .A2(new_n592), .ZN(G299));
  AND3_X1   g168(.A1(new_n530), .A2(KEYINPUT79), .A3(new_n532), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT79), .B1(new_n530), .B2(new_n532), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(G303));
  NAND2_X1  g171(.A1(new_n591), .A2(G87), .ZN(new_n597));
  INV_X1    g172(.A(G74), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n507), .B1(new_n520), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n540), .B2(G49), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(G288));
  NAND2_X1  g176(.A1(G73), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n520), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n523), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n540), .A2(G48), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(KEYINPUT81), .A3(new_n523), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G86), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n588), .B2(new_n590), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G305));
  NAND2_X1  g191(.A1(G72), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G60), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n520), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n523), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT82), .Z(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(G47), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n540), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G85), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n623), .C1(new_n624), .C2(new_n589), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n591), .A2(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n540), .A2(G54), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(new_n507), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n626), .B1(new_n634), .B2(G868), .ZN(G321));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NOR2_X1   g212(.A1(G168), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n581), .A2(new_n592), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT84), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(KEYINPUT84), .B2(new_n638), .ZN(G297));
  OAI21_X1  g218(.A(new_n642), .B1(KEYINPUT84), .B2(new_n638), .ZN(G280));
  INV_X1    g219(.A(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n634), .B1(new_n645), .B2(G860), .ZN(G148));
  OR3_X1    g221(.A1(new_n633), .A2(KEYINPUT85), .A3(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(KEYINPUT85), .B1(new_n633), .B2(G559), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G868), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g226(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g227(.A1(new_n488), .A2(new_n468), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n466), .A2(G135), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n478), .A2(G123), .ZN(new_n658));
  OR2_X1    g233(.A1(G99), .A2(G2105), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n659), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2096), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n662), .ZN(G156));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2435), .ZN(new_n665));
  XOR2_X1   g240(.A(G2427), .B(G2438), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT14), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT86), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(KEYINPUT86), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n676), .A2(G14), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G401));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2067), .B(G2678), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n681), .B1(new_n685), .B2(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2096), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n688), .A3(KEYINPUT17), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n687), .B(new_n691), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT87), .B(G2100), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT88), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n696), .A2(new_n697), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT20), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n699), .A2(new_n701), .A3(new_n704), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(G229));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G35), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G162), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT29), .B(G2090), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n715), .A2(G33), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n468), .A2(G103), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n466), .A2(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n723), .C1(new_n477), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n729), .A2(new_n715), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G160), .B2(new_n715), .ZN(new_n732));
  OR2_X1    g307(.A1(G29), .A2(G32), .ZN(new_n733));
  AOI22_X1  g308(.A1(G129), .A2(new_n478), .B1(new_n466), .B2(G141), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n468), .A2(G105), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(new_n715), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n728), .B1(new_n732), .B2(G2084), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n726), .B2(new_n727), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n715), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n715), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n745), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G21), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G168), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT92), .B(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n749), .A2(new_n750), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT93), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n661), .B2(new_n715), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n756), .B1(new_n769), .B2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n732), .A2(G2084), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n770), .B(new_n771), .C1(KEYINPUT95), .C2(new_n769), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n715), .A2(G26), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n466), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n478), .A2(G128), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n715), .ZN(new_n782));
  MUX2_X1   g357(.A(new_n775), .B(new_n782), .S(KEYINPUT28), .Z(new_n783));
  INV_X1    g358(.A(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n565), .A2(new_n746), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n746), .B2(G19), .ZN(new_n787));
  INV_X1    g362(.A(G1341), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n746), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n634), .B2(new_n746), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1348), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT97), .B(G1956), .Z(new_n794));
  OAI21_X1  g369(.A(KEYINPUT23), .B1(new_n640), .B2(new_n746), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n746), .A2(G20), .ZN(new_n796));
  MUX2_X1   g371(.A(KEYINPUT23), .B(new_n795), .S(new_n796), .Z(new_n797));
  OAI211_X1 g372(.A(new_n790), .B(new_n793), .C1(new_n794), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n794), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n772), .A2(new_n773), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n774), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G23), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n802), .A2(G16), .A3(G23), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n803), .B(new_n804), .C1(G288), .C2(new_n746), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT33), .B(G1976), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n746), .A2(G6), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n615), .B2(new_n746), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G22), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G166), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n715), .A2(G25), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n466), .A2(G131), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G119), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(new_n715), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  MUX2_X1   g406(.A(G24), .B(G290), .S(G16), .Z(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(G1986), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G1986), .B2(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n820), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n820), .A2(KEYINPUT91), .A3(new_n830), .A4(new_n834), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n819), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g416(.A(KEYINPUT36), .B(new_n819), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n719), .B(new_n801), .C1(new_n841), .C2(new_n842), .ZN(G150));
  INV_X1    g418(.A(G150), .ZN(G311));
  AOI22_X1  g419(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n512), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n548), .A2(G93), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT98), .B(G55), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n540), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n634), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n560), .B(KEYINPUT75), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n850), .B1(new_n855), .B2(new_n555), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n850), .B(new_n555), .C1(new_n561), .C2(new_n563), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT39), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n854), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n852), .B1(new_n861), .B2(G860), .ZN(G145));
  XOR2_X1   g437(.A(new_n474), .B(new_n661), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n738), .B(KEYINPUT99), .Z(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(new_n505), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n505), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n780), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n781), .A3(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n725), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(KEYINPUT100), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n477), .A2(G118), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n467), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .C1(G106), .C2(G2105), .ZN(new_n878));
  AOI22_X1  g453(.A1(G130), .A2(new_n478), .B1(new_n466), .B2(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n654), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n827), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT103), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n869), .A2(new_n725), .A3(new_n870), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT101), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n874), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(new_n874), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n864), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  INV_X1    g467(.A(new_n864), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n872), .A2(new_n873), .B1(new_n885), .B2(new_n886), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n888), .B(new_n893), .C1(new_n882), .C2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g472(.A(new_n649), .B(new_n859), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n640), .A2(new_n633), .ZN(new_n899));
  NAND4_X1  g474(.A1(G299), .A2(new_n630), .A3(new_n629), .A4(new_n632), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT104), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT41), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n898), .A2(new_n909), .A3(new_n901), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n615), .B(G166), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G288), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n919), .B2(KEYINPUT105), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(KEYINPUT105), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n917), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  INV_X1    g498(.A(new_n914), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n903), .A2(new_n908), .A3(new_n924), .A4(new_n910), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n915), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n915), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n850), .A2(new_n637), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(G171), .A2(KEYINPUT107), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n856), .B2(new_n858), .ZN(new_n936));
  OAI21_X1  g511(.A(G286), .B1(KEYINPUT107), .B2(G171), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n850), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n564), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n857), .A3(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n940), .A2(new_n857), .A3(new_n934), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n934), .B1(new_n940), .B2(new_n857), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n945), .C1(new_n904), .C2(new_n905), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n943), .A2(new_n944), .A3(new_n937), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n936), .B2(new_n941), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n901), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n933), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n942), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT108), .B1(new_n951), .B2(new_n901), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n922), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n922), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(KEYINPUT109), .A3(new_n922), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n932), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(KEYINPUT108), .ZN(new_n964));
  INV_X1    g539(.A(new_n952), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n954), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n922), .B1(new_n950), .B2(new_n952), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n892), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n955), .A2(new_n961), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT110), .B1(new_n973), .B2(new_n932), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n975), .B(KEYINPUT44), .C1(new_n970), .C2(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n974), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(KEYINPUT127), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n505), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT111), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT112), .B(G40), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n469), .A2(new_n473), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n738), .B(G1996), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n780), .B(new_n784), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n826), .A2(new_n829), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n826), .A2(new_n829), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(G1986), .B2(G290), .ZN(new_n998));
  OR2_X1    g573(.A1(G290), .A2(G1986), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n980), .A2(KEYINPUT113), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n491), .B2(new_n504), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT116), .B(new_n988), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n982), .B(G1384), .C1(new_n491), .C2(new_n504), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(G2078), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n505), .B2(new_n979), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT113), .B(G1384), .C1(new_n491), .C2(new_n504), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n988), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n988), .A2(KEYINPUT45), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1006), .A2(new_n1009), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n987), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n750), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT124), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n980), .A2(new_n982), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n754), .A3(new_n988), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT125), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1008), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1027), .B2(new_n1008), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1016), .A2(KEYINPUT124), .A3(new_n1021), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1006), .A2(new_n1026), .A3(new_n1015), .ZN(new_n1036));
  INV_X1    g611(.A(new_n759), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1020), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT117), .B(G2084), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT51), .B(G8), .C1(new_n1042), .C2(G286), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G168), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1036), .A2(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1044), .B(new_n1047), .C1(new_n1048), .C2(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1035), .B1(new_n1052), .B2(KEYINPUT62), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  NAND4_X1  g629(.A1(G303), .A2(new_n1054), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT79), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n548), .A2(G88), .B1(new_n523), .B2(new_n522), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n531), .B1(new_n1057), .B2(new_n514), .ZN(new_n1058));
  INV_X1    g633(.A(new_n532), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n530), .A2(KEYINPUT79), .A3(new_n532), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(KEYINPUT55), .A3(G8), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT114), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(G8), .A3(new_n1061), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1055), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1055), .A2(new_n1063), .A3(KEYINPUT115), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1025), .A2(new_n988), .A3(new_n1026), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n815), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1020), .B2(G2090), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1045), .B1(new_n1005), .B2(new_n988), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n548), .A2(G86), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G1981), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n612), .A2(G1981), .A3(new_n614), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n612), .A2(G1981), .A3(new_n614), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1081), .A3(KEYINPUT49), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n918), .A2(G1976), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1077), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1012), .A3(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT52), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1087), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1001), .A2(KEYINPUT50), .A3(new_n1004), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n987), .B1(new_n1002), .B2(new_n1017), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1045), .B1(new_n1098), .B2(new_n1073), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1076), .B(new_n1094), .C1(new_n1099), .C2(new_n1067), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1043), .A2(new_n1049), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT56), .B(G2072), .Z(new_n1105));
  NOR4_X1   g680(.A1(new_n1104), .A2(new_n1007), .A3(new_n987), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n591), .A2(G91), .ZN(new_n1110));
  INV_X1    g685(.A(new_n586), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n577), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT57), .B(new_n592), .C1(new_n578), .C2(new_n580), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(KEYINPUT119), .A3(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1109), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1005), .A2(new_n784), .A3(new_n988), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1348), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(new_n633), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1109), .A2(new_n1119), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1120), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n988), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(KEYINPUT50), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1130), .A2(G1956), .B1(new_n1072), .B2(new_n1105), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1117), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1115), .B(KEYINPUT57), .C1(new_n592), .C2(new_n577), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT119), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1109), .A2(KEYINPUT122), .A3(new_n1137), .A4(new_n1119), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1138), .A3(KEYINPUT61), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1072), .A2(G1996), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT58), .B(G1341), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1005), .B2(new_n988), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n565), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT121), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1145), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n565), .B(new_n1147), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1122), .A2(new_n1123), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n633), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1109), .A2(KEYINPUT122), .A3(new_n1154), .A4(new_n1119), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1151), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n634), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1153), .B(new_n1155), .C1(new_n1157), .C2(new_n1152), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1127), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1074), .A2(G8), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1067), .A2(new_n1099), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1087), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n983), .A2(G40), .A3(G160), .A4(new_n1009), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1021), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  OAI211_X1 g742(.A(KEYINPUT54), .B(new_n1167), .C1(new_n1034), .C2(G171), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1159), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1166), .A2(G171), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1033), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT124), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1031), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1173), .B2(G301), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1174), .A2(new_n1175), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1053), .A2(new_n1103), .B1(new_n1169), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1042), .A2(G8), .A3(G168), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1094), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT63), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1087), .A2(new_n1089), .A3(new_n918), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1085), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1077), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1055), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1099), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1045), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(G168), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1163), .B1(new_n1190), .B2(new_n1076), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1178), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(new_n1067), .B2(new_n1099), .ZN(new_n1194));
  NOR4_X1   g769(.A1(new_n1194), .A2(new_n1048), .A3(new_n1045), .A4(G286), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1094), .B1(new_n1195), .B2(new_n1161), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1184), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1163), .B1(new_n1186), .B2(new_n1160), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1198), .A2(G168), .A3(new_n1189), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1197), .B1(new_n1199), .B2(KEYINPUT63), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1196), .A2(new_n1200), .A3(KEYINPUT118), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1192), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1000), .B1(new_n1177), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n989), .A2(G1996), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1205));
  INV_X1    g780(.A(new_n989), .ZN(new_n1206));
  INV_X1    g781(.A(new_n991), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1206), .B1(new_n738), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT47), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n989), .A2(new_n999), .ZN(new_n1212));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1206), .A2(new_n997), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g791(.A1(new_n993), .A2(new_n995), .B1(new_n784), .B2(new_n781), .ZN(new_n1217));
  OR2_X1    g792(.A1(new_n1217), .A2(new_n989), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1211), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n978), .B1(new_n1203), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1000), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1164), .B1(new_n1052), .B2(KEYINPUT62), .ZN(new_n1222));
  OAI211_X1 g797(.A(G171), .B(new_n1034), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1052), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1159), .A2(new_n1168), .A3(new_n1164), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1222), .A2(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1192), .A2(new_n1201), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1221), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1219), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1229), .A2(KEYINPUT127), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1220), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g807(.A1(G229), .A2(new_n461), .ZN(new_n1234));
  NOR2_X1   g808(.A1(G401), .A2(G227), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n896), .A2(new_n973), .A3(new_n1234), .A4(new_n1235), .ZN(G225));
  INV_X1    g810(.A(G225), .ZN(G308));
endmodule


