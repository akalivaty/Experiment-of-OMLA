//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NOR2_X1   g0043(.A1(G20), .A2(G33), .ZN(new_n244));
  AOI22_X1  g0044(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n207), .A2(G33), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n207), .A3(G1), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n250), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n207), .A2(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n202), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n254), .A2(new_n256), .B1(new_n202), .B2(new_n253), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT71), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n251), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(KEYINPUT9), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1698), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n267), .A2(G222), .B1(new_n270), .B2(G77), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n265), .B2(new_n266), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G41), .A2(G45), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n213), .B1(new_n285), .B2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT65), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n277), .A2(new_n288), .A3(new_n280), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n283), .B1(new_n290), .B2(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n279), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g0092(.A(KEYINPUT70), .B(G200), .Z(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n262), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT72), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n279), .A2(new_n291), .A3(new_n299), .A4(G190), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(new_n261), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n260), .B1(new_n251), .B2(new_n257), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n296), .A2(new_n301), .A3(new_n302), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n298), .A3(new_n300), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n262), .A2(new_n295), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n292), .A2(G169), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n292), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n258), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n249), .A2(new_n213), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n252), .A2(G1), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G77), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n255), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n319), .A2(new_n322), .B1(G77), .B2(new_n318), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  INV_X1    g0124(.A(new_n244), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n247), .A2(new_n325), .B1(new_n207), .B2(new_n320), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT15), .B(G87), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT68), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n246), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n331), .B2(new_n316), .ZN(new_n332));
  INV_X1    g0132(.A(new_n326), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n327), .A2(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n327), .A2(KEYINPUT68), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(new_n246), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n323), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G244), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n287), .B2(new_n289), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT66), .B1(new_n341), .B2(new_n283), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n277), .A2(new_n288), .A3(new_n280), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n288), .B1(new_n277), .B2(new_n280), .ZN(new_n344));
  OAI21_X1  g0144(.A(G244), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT66), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n282), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n273), .A2(G238), .B1(new_n270), .B2(G107), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n270), .A2(KEYINPUT67), .A3(new_n231), .A4(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT67), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n267), .B2(G232), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n278), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n294), .B1(new_n348), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n339), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(G169), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n348), .A2(G179), .A3(new_n354), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n339), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n311), .A2(new_n315), .A3(new_n358), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G68), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n317), .A2(G20), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n244), .A2(G50), .B1(G20), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n320), .B2(new_n246), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT11), .A3(new_n250), .ZN(new_n369));
  INV_X1    g0169(.A(new_n255), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n254), .A2(G68), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT11), .B1(new_n368), .B2(new_n250), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(KEYINPUT14), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n343), .A2(new_n344), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT73), .B1(new_n287), .B2(new_n289), .ZN(new_n382));
  OAI21_X1  g0182(.A(G238), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(G226), .B(new_n272), .C1(new_n268), .C2(new_n269), .ZN(new_n384));
  OAI211_X1 g0184(.A(G232), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n283), .B1(new_n387), .B2(new_n278), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n379), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G238), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n380), .B1(new_n343), .B2(new_n344), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n289), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n387), .A2(new_n278), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n282), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT13), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n377), .B(new_n378), .C1(new_n389), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n383), .A2(new_n379), .A3(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n393), .B2(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n399), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n378), .B1(new_n402), .B2(new_n377), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT75), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n378), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n389), .A2(new_n396), .ZN(new_n406));
  INV_X1    g0206(.A(new_n377), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n397), .A4(new_n400), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n374), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n402), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G190), .B2(new_n402), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n374), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n247), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n370), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(KEYINPUT77), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n319), .B1(new_n418), .B2(KEYINPUT77), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n419), .A2(new_n420), .B1(new_n253), .B2(new_n247), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G58), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n364), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n424), .B2(new_n201), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n244), .A2(G159), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n268), .A2(new_n269), .A3(G20), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .A3(KEYINPUT7), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n265), .A2(new_n207), .A3(new_n266), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n266), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n427), .B1(new_n436), .B2(G68), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n316), .B1(new_n437), .B2(KEYINPUT16), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n431), .A2(new_n432), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n364), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n441), .B2(new_n427), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n422), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G223), .B(new_n272), .C1(new_n268), .C2(new_n269), .ZN(new_n444));
  OAI211_X1 g0244(.A(G226), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n445));
  INV_X1    g0245(.A(G87), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(new_n445), .C1(new_n264), .C2(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n447), .A2(new_n278), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n282), .B1(new_n286), .B2(new_n231), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n375), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n447), .B2(new_n278), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n313), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT18), .B1(new_n443), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n427), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n434), .A2(new_n430), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT76), .B1(new_n428), .B2(KEYINPUT7), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n434), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT16), .B(new_n455), .C1(new_n458), .C2(new_n364), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n250), .A3(new_n442), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n421), .ZN(new_n461));
  INV_X1    g0261(.A(new_n453), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n451), .A2(new_n297), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G200), .B2(new_n451), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n466), .A3(new_n421), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n460), .A2(new_n466), .A3(KEYINPUT17), .A4(new_n421), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n454), .A2(new_n464), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NOR4_X1   g0271(.A1(new_n363), .A2(new_n411), .A3(new_n416), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n318), .B1(new_n334), .B2(new_n335), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n207), .B1(new_n386), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G87), .A2(G97), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n475), .A2(new_n478), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n265), .A2(new_n266), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n207), .A3(G68), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n316), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n206), .A2(G33), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n316), .A2(new_n318), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n329), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(G250), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n206), .B2(G45), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n277), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n277), .A3(new_n490), .ZN(new_n495));
  INV_X1    g0295(.A(G45), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G1), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n494), .A2(new_n495), .B1(G274), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n264), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n267), .A2(KEYINPUT81), .A3(G238), .ZN(new_n504));
  OAI211_X1 g0304(.A(G238), .B(new_n272), .C1(new_n268), .C2(new_n269), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n498), .B(new_n313), .C1(new_n508), .C2(new_n277), .ZN(new_n509));
  INV_X1    g0309(.A(new_n495), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n206), .A2(G45), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n493), .B1(new_n281), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n503), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT81), .B1(new_n267), .B2(G238), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n505), .A2(new_n506), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n516), .B2(new_n278), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n489), .B(new_n509), .C1(new_n517), .C2(G169), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n498), .B(G190), .C1(new_n508), .C2(new_n277), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n486), .A2(new_n446), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n473), .A2(new_n483), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n521), .C1(new_n517), .C2(new_n293), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n477), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  XNOR2_X1  g0325(.A(G97), .B(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n528), .A2(new_n207), .B1(new_n320), .B2(new_n325), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n477), .B1(new_n440), .B2(new_n434), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n250), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n318), .A2(G97), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n487), .B2(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(G244), .C1(new_n269), .C2(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n340), .B1(new_n265), .B2(new_n266), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(KEYINPUT4), .ZN(new_n540));
  OAI21_X1  g0340(.A(G250), .B1(new_n268), .B2(new_n269), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n272), .B1(new_n541), .B2(KEYINPUT4), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n278), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(KEYINPUT5), .A2(G41), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n497), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(G257), .A3(new_n277), .ZN(new_n548));
  OR2_X1    g0348(.A1(KEYINPUT5), .A2(G41), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n511), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G274), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT78), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n543), .A2(new_n553), .A3(new_n313), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n534), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n552), .ZN(new_n558));
  AOI21_X1  g0358(.A(G169), .B1(new_n543), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n524), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(KEYINPUT79), .A3(new_n534), .A4(new_n556), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n543), .A2(new_n553), .A3(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n531), .A2(new_n533), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n543), .A2(G190), .A3(new_n558), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n523), .A2(new_n560), .A3(new_n562), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT20), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n207), .A2(new_n500), .ZN(new_n570));
  INV_X1    g0370(.A(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n538), .B1(new_n571), .B2(G33), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(new_n207), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n569), .B1(new_n573), .B2(new_n316), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n264), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(G20), .B1(new_n575), .B2(new_n538), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT20), .B(new_n250), .C1(new_n576), .C2(new_n570), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n486), .A2(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n318), .A2(new_n500), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n375), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n272), .C1(new_n268), .C2(new_n269), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n584));
  OAI211_X1 g0384(.A(G264), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(KEYINPUT82), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT82), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n273), .B2(G264), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n278), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n550), .A2(new_n278), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G270), .B1(G274), .B2(new_n550), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT21), .B1(new_n582), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n592), .A2(G190), .ZN(new_n595));
  AOI21_X1  g0395(.A(G200), .B1(new_n589), .B2(new_n591), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n578), .B(new_n581), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n578), .A2(new_n581), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(new_n598), .A3(KEYINPUT21), .A4(G169), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(G179), .A3(new_n589), .A4(new_n591), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(KEYINPUT83), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT83), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n594), .B(new_n597), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n207), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n477), .A2(KEYINPUT23), .A3(G20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n501), .A2(new_n207), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n207), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT22), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT22), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n481), .A2(new_n612), .A3(new_n207), .A4(G87), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(KEYINPUT24), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n316), .B1(new_n614), .B2(KEYINPUT24), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n317), .A2(G20), .A3(new_n477), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT25), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(G107), .B2(new_n487), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G294), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n541), .C2(G1698), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n278), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n590), .A2(G264), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n551), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(G179), .A3(new_n551), .A4(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n627), .A2(new_n412), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n627), .A2(G190), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n617), .B(new_n620), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n568), .A2(new_n603), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n472), .A2(new_n636), .ZN(G372));
  NOR3_X1   g0437(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n374), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n407), .B1(new_n398), .B2(new_n399), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n378), .B1(new_n406), .B2(G179), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n409), .B1(new_n644), .B2(new_n408), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n401), .A2(KEYINPUT75), .A3(new_n403), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n362), .B1(new_n414), .B2(new_n374), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n469), .A2(new_n470), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n641), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n311), .ZN(new_n653));
  OAI211_X1 g0453(.A(KEYINPUT84), .B(new_n315), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT84), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n651), .B1(new_n411), .B2(new_n648), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n653), .B1(new_n656), .B2(new_n640), .ZN(new_n657));
  INV_X1    g0457(.A(new_n315), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n634), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n617), .A2(new_n620), .B1(new_n628), .B2(new_n629), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n599), .A2(new_n600), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n662), .A2(new_n663), .A3(new_n593), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n568), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n557), .A2(new_n559), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n523), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n518), .A2(new_n522), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n560), .B2(new_n562), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n668), .B(new_n518), .C1(new_n670), .C2(new_n666), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n472), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(new_n317), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .A3(G20), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT27), .B1(new_n674), .B2(G20), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n598), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n663), .A2(new_n593), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n603), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n679), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n631), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT86), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n617), .B2(new_n620), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT85), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n631), .A3(new_n634), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(KEYINPUT86), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n686), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n683), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n594), .B1(new_n601), .B2(new_n602), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n684), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n693), .A2(new_n696), .B1(new_n662), .B2(new_n684), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n210), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n206), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n476), .A2(new_n477), .A3(new_n500), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(new_n703), .B1(new_n217), .B2(new_n700), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  NOR2_X1   g0505(.A1(new_n592), .A2(new_n313), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n625), .A2(new_n626), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n543), .A2(new_n558), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n707), .A3(new_n709), .A4(new_n517), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  INV_X1    g0511(.A(new_n517), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(new_n627), .A3(new_n563), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n592), .A2(new_n313), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n710), .A2(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n710), .A2(new_n711), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n679), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n679), .C1(new_n715), .C2(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n560), .A2(new_n562), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n567), .A2(new_n518), .A3(new_n522), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n722), .A2(new_n635), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n603), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(new_n684), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT87), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n636), .A2(KEYINPUT87), .A3(new_n684), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n721), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n684), .B1(new_n665), .B2(new_n671), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n594), .B(new_n631), .C1(new_n601), .C2(new_n602), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n560), .A2(new_n562), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n567), .A2(new_n518), .A3(new_n522), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n634), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n722), .A2(new_n666), .A3(new_n523), .ZN(new_n740));
  INV_X1    g0540(.A(new_n518), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n534), .A2(new_n556), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n518), .A3(new_n522), .A4(new_n561), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(KEYINPUT26), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT88), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n740), .A2(new_n744), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n679), .B1(new_n749), .B2(new_n739), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n732), .B1(new_n735), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n705), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n682), .A2(G330), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n252), .A2(G20), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT89), .Z(new_n758));
  NAND2_X1  g0558(.A1(new_n701), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n683), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n213), .B1(G20), .B2(new_n375), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n313), .A2(new_n412), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n481), .B1(new_n766), .B2(new_n364), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n294), .A2(new_n313), .ZN(new_n768));
  INV_X1    g0568(.A(new_n765), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n477), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n207), .B1(new_n773), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n767), .B(new_n772), .C1(G97), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n297), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n768), .A2(KEYINPUT93), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT93), .B1(new_n768), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G87), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n313), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT90), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n765), .A2(new_n773), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(KEYINPUT32), .A3(G159), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n786), .A2(G58), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n777), .A2(new_n764), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT92), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(KEYINPUT92), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n765), .A2(new_n784), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G50), .A2(new_n799), .B1(new_n806), .B2(G77), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n776), .A2(new_n783), .A3(new_n793), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n782), .A2(G303), .ZN(new_n809));
  INV_X1    g0609(.A(new_n766), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT33), .B(G317), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT94), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n813), .A2(new_n814), .B1(new_n815), .B2(new_n785), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n481), .B1(new_n791), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n774), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n806), .B2(G311), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n799), .A2(G326), .B1(new_n770), .B2(G283), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n809), .A2(new_n817), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n763), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G13), .A2(G33), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n762), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n699), .A2(new_n270), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G355), .B1(new_n500), .B2(new_n699), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n217), .A2(G45), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n242), .B2(G45), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n699), .A2(new_n481), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n759), .B(new_n824), .C1(new_n828), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  INV_X1    g0637(.A(new_n827), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n682), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n761), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n762), .A2(new_n825), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G303), .A2(new_n799), .B1(new_n806), .B2(G116), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n270), .B1(new_n788), .B2(new_n845), .C1(new_n785), .C2(new_n819), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G97), .B2(new_n775), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n810), .A2(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n810), .A2(KEYINPUT97), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(G283), .B1(new_n770), .B2(G87), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n844), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G107), .B2(new_n782), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n786), .A2(G143), .B1(G150), .B2(new_n810), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n855), .B2(new_n798), .C1(new_n789), .C2(new_n805), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n481), .B1(new_n788), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT98), .Z(new_n861));
  AOI22_X1  g0661(.A1(new_n770), .A2(G68), .B1(G58), .B2(new_n775), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(new_n781), .C2(new_n202), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n856), .B2(new_n857), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n853), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n760), .B1(G77), .B2(new_n843), .C1(new_n865), .C2(new_n763), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n679), .B(new_n339), .C1(new_n359), .C2(new_n360), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n339), .A2(new_n684), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n358), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(new_n362), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n866), .B1(new_n825), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n733), .B(new_n870), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n732), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n760), .B1(new_n732), .B2(new_n873), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G384));
  INV_X1    g0677(.A(new_n528), .ZN(new_n878));
  OAI211_X1 g0678(.A(G116), .B(new_n214), .C1(new_n878), .C2(KEYINPUT35), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(KEYINPUT35), .B2(new_n878), .ZN(new_n880));
  XNOR2_X1  g0680(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  OR3_X1    g0682(.A1(new_n216), .A2(new_n320), .A3(new_n424), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n202), .A2(G68), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n206), .B(G13), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n374), .A2(new_n684), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n647), .A2(new_n415), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n411), .B2(new_n416), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n871), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n721), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT87), .B1(new_n636), .B2(new_n684), .ZN(new_n893));
  AND4_X1   g0693(.A1(KEYINPUT87), .A2(new_n724), .A3(new_n725), .A4(new_n684), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n455), .B1(new_n458), .B2(new_n364), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n439), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n422), .B1(new_n438), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n677), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n640), .B2(new_n651), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n461), .A2(new_n462), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n677), .B(KEYINPUT100), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n461), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n467), .ZN(new_n907));
  INV_X1    g0707(.A(new_n677), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n450), .B2(new_n452), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n467), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n896), .B1(new_n902), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n471), .A2(new_n900), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n911), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n891), .A2(new_n895), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n903), .A2(new_n905), .A3(new_n467), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  INV_X1    g0722(.A(new_n905), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n907), .B1(new_n471), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n895), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n895), .A2(new_n472), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n927), .B(new_n928), .Z(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n731), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT88), .B1(new_n750), .B2(KEYINPUT29), .ZN(new_n931));
  AND4_X1   g0731(.A1(KEYINPUT88), .A2(new_n745), .A3(KEYINPUT29), .A4(new_n684), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n472), .B(new_n735), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT101), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT101), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n752), .A2(new_n935), .A3(new_n472), .A4(new_n735), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n660), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n889), .A2(new_n890), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n684), .B(new_n870), .C1(new_n665), .C2(new_n671), .ZN(new_n939));
  INV_X1    g0739(.A(new_n867), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n917), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n640), .A2(new_n904), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n647), .A2(new_n679), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n914), .B2(new_n915), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT39), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n916), .B(new_n950), .C1(new_n924), .C2(KEYINPUT38), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n946), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n937), .B(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n930), .A2(new_n954), .B1(new_n206), .B2(new_n756), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n930), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n886), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT102), .ZN(G367));
  NOR2_X1   g0758(.A1(new_n684), .A2(new_n521), .ZN(new_n959));
  MUX2_X1   g0759(.A(new_n523), .B(new_n741), .S(new_n959), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n838), .ZN(new_n961));
  INV_X1    g0761(.A(new_n828), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n833), .B2(new_n235), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n329), .A2(new_n699), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n759), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(G143), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n798), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n771), .A2(new_n320), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G159), .C2(new_n850), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n481), .B1(new_n788), .B2(new_n855), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n806), .B2(G50), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n782), .A2(G58), .ZN(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n785), .A2(new_n973), .B1(new_n774), .B2(new_n364), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT109), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n781), .A2(new_n977), .A3(new_n500), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n771), .A2(new_n571), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G294), .B2(new_n850), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n781), .B2(new_n500), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n481), .B1(new_n791), .B2(G317), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n477), .B2(new_n774), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n799), .B2(G311), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n806), .A2(G283), .B1(G303), .B2(new_n786), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n976), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT47), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n762), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n965), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n961), .B1(new_n991), .B2(KEYINPUT110), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT110), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n758), .A2(G1), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n696), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n631), .B2(new_n679), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n667), .A2(new_n679), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT104), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n534), .A2(new_n679), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n737), .A2(new_n567), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT103), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(KEYINPUT103), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n996), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1000), .B(KEYINPUT103), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n998), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT45), .B1(new_n1008), .B2(new_n697), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT106), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1008), .A2(new_n697), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1013), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n996), .B2(new_n1003), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1014), .A2(new_n1016), .B1(KEYINPUT106), .B2(KEYINPUT44), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1010), .B(new_n1017), .C1(KEYINPUT107), .C2(new_n694), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1013), .B1(new_n1008), .B2(new_n697), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n996), .A2(new_n1003), .A3(new_n1015), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n693), .A2(new_n696), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT108), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n995), .C1(new_n1026), .C2(new_n683), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n683), .A2(new_n1026), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  NAND4_X1  g0829(.A1(new_n1018), .A2(new_n1024), .A3(new_n753), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n753), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n700), .B(KEYINPUT41), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n994), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1003), .A2(new_n995), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT42), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n1008), .A2(new_n662), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n679), .B1(new_n1037), .B2(new_n737), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n694), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1008), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT105), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1039), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n1045), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n993), .B1(new_n1034), .B2(new_n1053), .ZN(G387));
  OR2_X1    g0854(.A1(new_n1029), .A2(new_n753), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1029), .A2(new_n753), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n700), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n693), .A2(new_n838), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n829), .A2(new_n702), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(G107), .B2(new_n210), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n232), .A2(G45), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n417), .A2(new_n202), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT112), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT111), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n496), .B1(new_n364), .B2(new_n320), .C1(new_n702), .C2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n702), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n834), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1060), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n760), .B1(new_n1069), .B2(new_n962), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT113), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n481), .B1(new_n791), .B2(G326), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n850), .A2(G311), .B1(G317), .B2(new_n786), .ZN(new_n1073));
  INV_X1    g0873(.A(G303), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n805), .C1(new_n815), .C2(new_n798), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n782), .A2(G294), .B1(G283), .B2(new_n775), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1072), .B1(new_n500), .B2(new_n771), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n270), .B(new_n979), .C1(G150), .C2(new_n791), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n782), .A2(G77), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT114), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n799), .A2(G159), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n806), .A2(G68), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n785), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G50), .A2(new_n1090), .B1(new_n810), .B2(new_n417), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n329), .A2(new_n775), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1082), .A2(new_n1083), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1058), .B(new_n1071), .C1(new_n762), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1029), .B2(new_n994), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1057), .A2(new_n1096), .ZN(G393));
  NAND3_X1  g0897(.A1(new_n1010), .A2(new_n1017), .A3(new_n1040), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n694), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n994), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n833), .A2(new_n239), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n962), .B1(G97), .B2(new_n699), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n759), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n481), .B(new_n772), .C1(G322), .C2(new_n791), .ZN(new_n1106));
  INV_X1    g0906(.A(G283), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n781), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT115), .Z(new_n1109));
  INV_X1    g0909(.A(new_n850), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1110), .A2(new_n1074), .B1(new_n500), .B2(new_n774), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n799), .A2(G317), .B1(G311), .B2(new_n1090), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(G294), .C2(new_n806), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n798), .A2(new_n973), .B1(new_n789), .B2(new_n785), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n481), .B1(new_n774), .B2(new_n320), .C1(new_n966), .C2(new_n788), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n770), .B2(G87), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n247), .B2(new_n805), .C1(new_n1110), .C2(new_n202), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G68), .B2(new_n782), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1109), .A2(new_n1114), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1105), .B1(new_n1008), .B2(new_n838), .C1(new_n763), .C2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1101), .A2(new_n1102), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1098), .A2(new_n1099), .B1(G1), .B2(new_n758), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1122), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1056), .A2(new_n1099), .A3(new_n1098), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1030), .A2(new_n1128), .A3(new_n700), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT117), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT117), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1030), .A2(new_n1128), .A3(new_n1131), .A4(new_n700), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n945), .B1(new_n938), .B2(new_n941), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n949), .A2(new_n951), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n869), .A2(new_n362), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n750), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1137), .A2(new_n940), .B1(new_n889), .B2(new_n890), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n946), .A2(new_n925), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1134), .A2(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n891), .A2(G330), .A3(new_n895), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n889), .A2(new_n890), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n867), .B1(new_n750), .B2(new_n1136), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n946), .B(new_n925), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n1141), .C1(new_n1135), .C2(new_n1134), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n994), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n760), .B1(new_n417), .B2(new_n843), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n270), .B1(new_n788), .B2(new_n819), .C1(new_n785), .C2(new_n500), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G77), .B2(new_n775), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n806), .A2(G97), .B1(new_n770), .B2(G68), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n799), .A2(G283), .B1(new_n850), .B2(G107), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n783), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n782), .A2(G150), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n774), .A2(new_n789), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1110), .A2(new_n855), .B1(new_n771), .B2(new_n202), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n481), .B1(new_n788), .B2(new_n1161), .C1(new_n785), .C2(new_n859), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n798), .A2(new_n1163), .B1(new_n805), .B2(new_n1164), .ZN(new_n1165));
  OR4_X1    g0965(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1156), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1151), .B1(new_n1167), .B2(new_n762), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1135), .B2(new_n826), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1145), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n730), .A2(new_n731), .A3(new_n871), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1141), .B(new_n1170), .C1(new_n1171), .C2(new_n938), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n895), .A2(G330), .A3(new_n870), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n1144), .B1(new_n732), .B2(new_n891), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1174), .B2(new_n941), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n928), .A2(G330), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n934), .A2(new_n660), .A3(new_n936), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1149), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n700), .B1(new_n1178), .B2(new_n1149), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1150), .B(new_n1169), .C1(new_n1180), .C2(new_n1181), .ZN(G378));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n311), .A2(new_n315), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n677), .B1(new_n259), .B2(new_n261), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1183), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n944), .B2(new_n952), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n951), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n950), .B1(new_n913), .B2(new_n916), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n945), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n943), .A3(new_n1198), .A4(new_n942), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n920), .A2(new_n926), .A3(G330), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1194), .B(new_n1199), .C1(new_n927), .C2(new_n731), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AND4_X1   g1004(.A1(new_n660), .A2(new_n934), .A3(new_n936), .A4(new_n1176), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1148), .B2(new_n1175), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n700), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1198), .A2(new_n825), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n760), .B1(G50), .B2(new_n843), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1213));
  INV_X1    g1013(.A(G41), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n270), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n771), .A2(new_n423), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G116), .B2(new_n799), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n766), .A2(new_n571), .B1(new_n788), .B2(new_n1107), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1214), .B(new_n270), .C1(new_n785), .C2(new_n477), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G68), .C2(new_n775), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n806), .A2(new_n329), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1085), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n774), .A2(new_n973), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1163), .A2(new_n785), .B1(new_n766), .B2(new_n859), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n806), .C2(G137), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n1161), .B2(new_n798), .C1(new_n781), .C2(new_n1164), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n770), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1224), .B1(new_n1223), .B2(new_n1222), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1212), .B1(new_n1234), .B2(new_n762), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1204), .A2(new_n994), .B1(new_n1211), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1210), .A2(new_n1236), .ZN(G375));
  INV_X1    g1037(.A(new_n1178), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1033), .A3(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1172), .B(new_n994), .C1(new_n1174), .C2(new_n941), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT118), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1141), .B1(new_n1171), .B2(new_n938), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n940), .A3(new_n939), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT118), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n994), .A4(new_n1172), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n938), .A2(new_n826), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT119), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G107), .A2(new_n806), .B1(new_n850), .B2(G116), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1092), .C1(new_n819), .C2(new_n798), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n781), .A2(new_n571), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n270), .B1(new_n788), .B2(new_n1074), .C1(new_n785), .C2(new_n1107), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1250), .A2(new_n968), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n481), .B1(new_n774), .B2(new_n202), .C1(new_n1163), .C2(new_n788), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1254), .B(new_n1216), .C1(G150), .C2(new_n806), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n789), .B2(new_n781), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n786), .A2(G137), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n859), .B2(new_n798), .C1(new_n1110), .C2(new_n1164), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(KEYINPUT120), .B2(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1258), .A2(KEYINPUT120), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1253), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n763), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n759), .B(new_n1262), .C1(new_n364), .C2(new_n842), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1242), .A2(new_n1246), .B1(new_n1248), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1240), .A2(new_n1264), .ZN(G381));
  NAND3_X1  g1065(.A1(new_n1057), .A2(new_n840), .A3(new_n1096), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(G387), .A2(G384), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1264), .A4(new_n1240), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT121), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(G407));
  NAND2_X1  g1074(.A1(new_n678), .A2(G213), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G407), .A2(G213), .A3(new_n1277), .ZN(G409));
  AOI22_X1  g1078(.A1(new_n1123), .A2(new_n1126), .B1(new_n1129), .B2(KEYINPUT117), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G387), .A2(new_n1132), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1032), .B1(new_n1030), .B2(new_n753), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1049), .B(new_n1052), .C1(new_n1281), .C2(new_n994), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G390), .A2(new_n1282), .A3(new_n993), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n840), .B1(new_n1057), .B2(new_n1096), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1266), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1280), .A2(new_n1283), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G387), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1285), .A2(new_n1266), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(G390), .C1(new_n1289), .C2(KEYINPUT124), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1268), .A2(new_n1289), .A3(G387), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT60), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n700), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT60), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1248), .A2(new_n1263), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n876), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1296), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT60), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1302), .A2(new_n1238), .A3(new_n700), .A4(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(G384), .A3(new_n1264), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1210), .A2(G378), .A3(new_n1236), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1150), .A2(new_n1169), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1181), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1179), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1204), .A2(new_n1206), .A3(new_n1033), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1236), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n1276), .B(new_n1306), .C1(new_n1307), .C2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1307), .A2(new_n1313), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1306), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1275), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1317), .A2(new_n1321), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1275), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT123), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1301), .A2(new_n1305), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1276), .A2(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1325), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1319), .A2(new_n1324), .A3(new_n1327), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1323), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT61), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1293), .B1(new_n1322), .B2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1318), .A2(KEYINPUT63), .A3(new_n1275), .A4(new_n1319), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1331), .A2(new_n1332), .A3(new_n1335), .A4(new_n1292), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1320), .A2(KEYINPUT122), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT122), .B1(new_n1320), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT125), .B1(new_n1337), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT122), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1314), .B2(KEYINPUT63), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1320), .A2(KEYINPUT122), .A3(new_n1338), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT125), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1346), .A2(new_n1336), .A3(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1334), .B1(new_n1342), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(KEYINPUT127), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1334), .B(new_n1351), .C1(new_n1342), .C2(new_n1348), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(G405));
  XNOR2_X1  g1153(.A(new_n1292), .B(new_n1306), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(G375), .B(new_n1310), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1354), .B(new_n1355), .ZN(G402));
endmodule


