//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT75), .B1(new_n187), .B2(G128), .ZN(new_n188));
  AOI22_X1  g002(.A1(new_n188), .A2(KEYINPUT23), .B1(new_n187), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(KEYINPUT75), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT24), .B(G110), .Z(new_n195));
  OAI21_X1  g009(.A(KEYINPUT74), .B1(new_n190), .B2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n187), .A3(G128), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(new_n198), .A3(new_n191), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(new_n210), .B(G146), .C1(new_n205), .C2(new_n206), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n199), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n204), .A3(new_n208), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n211), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT73), .B(G902), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n218), .A3(new_n223), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n226), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n226), .B2(G234), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n225), .A2(new_n227), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n234), .A2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n241));
  INV_X1    g055(.A(G237), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n242), .A2(new_n221), .A3(G210), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n241), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G101), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n208), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n208), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n252), .B(new_n254), .C1(G128), .C2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT66), .A2(G131), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT66), .A2(G131), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G137), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .A3(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n261), .A2(G137), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n257), .A2(new_n258), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n262), .A2(new_n264), .A3(new_n274), .A4(new_n265), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n250), .A2(G146), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(new_n253), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT0), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n190), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT65), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n249), .A2(new_n251), .B1(KEYINPUT0), .B2(G128), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n285), .A4(new_n284), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n249), .A2(new_n251), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n279), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n270), .B1(new_n278), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n187), .A2(G116), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G119), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n187), .A2(KEYINPUT68), .A3(G116), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT68), .B1(new_n187), .B2(G116), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n299), .A3(G119), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n305), .A2(new_n306), .B1(G116), .B2(new_n187), .ZN(new_n307));
  INV_X1    g121(.A(new_n303), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n296), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n302), .A2(new_n303), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n308), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT28), .B1(new_n295), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n256), .A2(new_n266), .A3(new_n269), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n287), .A2(new_n293), .A3(new_n290), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n275), .A2(G131), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n266), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n311), .A2(KEYINPUT69), .A3(new_n312), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT69), .B1(new_n311), .B2(new_n312), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n307), .B(new_n303), .ZN(new_n328));
  INV_X1    g142(.A(new_n279), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n286), .A2(new_n255), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n292), .B1(new_n330), .B2(new_n289), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n331), .A3(new_n287), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n332), .B2(new_n270), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n247), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n328), .ZN(new_n336));
  OAI211_X1 g150(.A(KEYINPUT30), .B(new_n270), .C1(new_n278), .C2(new_n294), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n336), .B(new_n337), .C1(new_n321), .C2(KEYINPUT30), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT31), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n246), .B1(new_n321), .B2(new_n324), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(G472), .A2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT71), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT72), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT31), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n333), .B1(new_n315), .B2(new_n326), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(new_n247), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n353));
  INV_X1    g167(.A(new_n345), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n226), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n332), .A2(new_n270), .B1(new_n310), .B2(new_n313), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n315), .B2(new_n326), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n246), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n295), .A2(new_n314), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n295), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n316), .A2(new_n364), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n328), .B1(new_n366), .B2(new_n332), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n360), .B1(new_n368), .B2(new_n247), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n246), .B(new_n333), .C1(new_n315), .C2(new_n326), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G472), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n349), .A2(new_n350), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT32), .B(new_n354), .C1(new_n373), .C2(new_n335), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n240), .B1(new_n356), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G210), .B1(G237), .B2(G902), .ZN(new_n379));
  OAI211_X1 g193(.A(KEYINPUT5), .B(new_n297), .C1(new_n300), .C2(new_n301), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(G113), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G104), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(G107), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n384), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n386), .A2(G104), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n383), .A2(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n382), .A2(new_n312), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(G101), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n396), .A2(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n401), .B2(new_n328), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n402), .A2(KEYINPUT82), .A3(new_n404), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n294), .A2(G125), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(G125), .B2(new_n256), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G953), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n402), .A2(new_n404), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n395), .B(new_n403), .C1(new_n401), .C2(new_n328), .ZN(new_n418));
  AND4_X1   g232(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT6), .A4(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n402), .B2(new_n404), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n421), .B2(new_n418), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n410), .B(new_n415), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(new_n413), .B2(G953), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n418), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n382), .A2(new_n312), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n390), .A2(new_n393), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n395), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n403), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n412), .A2(new_n424), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n423), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n379), .B1(new_n436), .B2(KEYINPUT84), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n423), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n423), .A2(new_n435), .A3(new_n379), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n378), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G221), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT9), .B(G234), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G902), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n446), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G140), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n221), .A2(G227), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n396), .A2(G101), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n331), .A2(new_n455), .A3(new_n398), .A4(new_n287), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n250), .A2(KEYINPUT1), .A3(G146), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n291), .B2(new_n190), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n252), .A2(KEYINPUT78), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n255), .A2(new_n460), .A3(new_n248), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n394), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n429), .A2(new_n464), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n256), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n456), .A2(new_n465), .A3(new_n467), .A4(new_n278), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n463), .A2(new_n464), .B1(new_n466), .B2(new_n256), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n456), .A4(new_n278), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n463), .B1(new_n394), .B2(new_n256), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(new_n320), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n474), .B2(new_n320), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n453), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n278), .B1(new_n470), .B2(new_n456), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n452), .B(new_n480), .C1(new_n469), .C2(new_n472), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n449), .B1(new_n482), .B2(G469), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n473), .A2(new_n453), .A3(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n453), .B1(new_n473), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n448), .B(new_n226), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n447), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n383), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n202), .A2(new_n204), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G146), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n217), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n242), .A2(new_n221), .A3(G214), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G143), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G237), .A2(G953), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(G214), .C1(new_n496), .C2(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(KEYINPUT18), .A2(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT87), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(KEYINPUT87), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n500), .ZN(new_n506));
  INV_X1    g320(.A(new_n501), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT86), .B(new_n501), .C1(new_n498), .C2(new_n500), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n494), .B(new_n504), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n211), .A2(new_n210), .ZN(new_n511));
  AOI21_X1  g325(.A(G146), .B1(new_n205), .B2(new_n206), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n213), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n272), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n498), .A2(new_n500), .A3(new_n259), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n259), .B1(new_n498), .B2(new_n500), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n491), .B(new_n510), .C1(new_n514), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n491), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n494), .A2(new_n504), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n506), .A2(new_n507), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT86), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n506), .A2(new_n505), .A3(new_n507), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT19), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT19), .B1(new_n202), .B2(new_n204), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n208), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n498), .A2(new_n500), .A3(new_n259), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n531), .B(new_n211), .C1(new_n532), .C2(new_n519), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n523), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n489), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT20), .B(new_n539), .C1(new_n522), .C2(new_n535), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G475), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n510), .B1(new_n514), .B2(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n523), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n522), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n545), .B2(new_n446), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT88), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n522), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n516), .B(new_n259), .C1(new_n500), .C2(new_n498), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n532), .A2(new_n519), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n516), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n212), .A2(new_n214), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n491), .B1(new_n553), .B2(new_n510), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n446), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G475), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(new_n557), .C1(new_n538), .C2(new_n540), .ZN(new_n558));
  XNOR2_X1  g372(.A(G128), .B(G143), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n261), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT89), .ZN(new_n561));
  XOR2_X1   g375(.A(G116), .B(G122), .Z(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G107), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(KEYINPUT13), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n250), .A2(G128), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(G134), .C1(KEYINPUT13), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n559), .B(new_n261), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n299), .A2(KEYINPUT14), .A3(G122), .ZN(new_n569));
  OAI211_X1 g383(.A(G107), .B(new_n569), .C1(new_n562), .C2(KEYINPUT14), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n568), .B(new_n570), .C1(G107), .C2(new_n562), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n444), .A2(new_n233), .A3(G953), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n567), .B2(new_n571), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n226), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G478), .ZN(new_n577));
  NOR2_X1   g391(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n576), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n547), .A2(new_n558), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G234), .A2(G237), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n357), .A2(G953), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT21), .B(G898), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n221), .A2(G952), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n587), .A2(new_n588), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n376), .A2(new_n442), .A3(new_n488), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NOR2_X1   g407(.A1(new_n341), .A2(new_n342), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n327), .A2(new_n334), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n246), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n357), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT91), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(G472), .C1(new_n343), .C2(new_n357), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n346), .A2(new_n355), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n447), .ZN(new_n605));
  INV_X1    g419(.A(new_n240), .ZN(new_n606));
  INV_X1    g420(.A(new_n487), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n473), .A2(new_n478), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n452), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n473), .A2(new_n485), .A3(new_n453), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(G469), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n449), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT92), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n346), .A2(new_n355), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n599), .B2(new_n601), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n447), .B(new_n240), .C1(new_n483), .C2(new_n487), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT93), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n379), .B1(new_n423), .B2(new_n435), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n377), .B(new_n441), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n441), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(KEYINPUT94), .A3(new_n377), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n590), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n547), .A2(new_n558), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  INV_X1    g444(.A(new_n572), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(KEYINPUT95), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n574), .B2(new_n575), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n567), .A2(new_n571), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n631), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n573), .A3(new_n632), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n634), .A2(new_n637), .A3(G478), .A4(new_n226), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n576), .A2(new_n577), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT96), .B1(new_n629), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n643), .B(new_n640), .C1(new_n547), .C2(new_n558), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n622), .A2(new_n628), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  OAI21_X1  g462(.A(KEYINPUT97), .B1(new_n538), .B2(new_n540), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n491), .B1(new_n510), .B2(new_n533), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n528), .B1(new_n552), .B2(new_n551), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n491), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT20), .B1(new_n652), .B2(new_n539), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n536), .A2(new_n489), .A3(new_n537), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n582), .A2(new_n649), .A3(new_n656), .A4(new_n556), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n590), .B(new_n657), .C1(new_n627), .C2(new_n625), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n622), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  INV_X1    g475(.A(new_n234), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n230), .B2(new_n231), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n219), .B(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n238), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n584), .A2(new_n590), .A3(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n617), .A2(new_n442), .A3(new_n488), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  AND3_X1   g485(.A1(new_n649), .A2(new_n656), .A3(new_n556), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n589), .A2(new_n585), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT98), .B(G900), .Z(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n587), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n672), .A2(new_n673), .A3(new_n582), .A4(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT100), .B1(new_n657), .B2(new_n678), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n356), .A2(new_n375), .ZN(new_n683));
  INV_X1    g497(.A(new_n667), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n605), .B(new_n684), .C1(new_n607), .C2(new_n613), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n627), .A2(new_n625), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  NAND2_X1  g503(.A1(new_n440), .A2(new_n441), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n368), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n247), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n363), .A2(new_n358), .A3(new_n247), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(G902), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n598), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n345), .B1(new_n594), .B2(new_n596), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n698), .B2(KEYINPUT32), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n356), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n547), .A2(new_n558), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n583), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n377), .A3(new_n667), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n692), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n678), .B(new_n705), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n488), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n707), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n704), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT103), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  AOI211_X1 g530(.A(new_n678), .B(new_n640), .C1(new_n547), .C2(new_n558), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n686), .A2(new_n683), .A3(new_n687), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  OAI21_X1  g533(.A(new_n226), .B1(new_n484), .B2(new_n486), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n448), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n473), .A2(new_n485), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n452), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n473), .A2(new_n453), .A3(new_n478), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n722), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n226), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n723), .A2(new_n729), .A3(new_n605), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n729), .A3(new_n732), .A4(new_n605), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n628), .A3(new_n376), .A4(new_n645), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n376), .A3(new_n658), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AOI21_X1  g553(.A(new_n730), .B1(new_n625), .B2(new_n627), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n683), .A3(new_n668), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  OR2_X1    g556(.A1(new_n359), .A2(new_n247), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n345), .B1(new_n594), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n597), .B2(new_n598), .ZN(new_n746));
  OAI211_X1 g560(.A(KEYINPUT106), .B(G472), .C1(new_n343), .C2(new_n357), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n235), .A2(new_n749), .A3(new_n239), .ZN(new_n750));
  INV_X1    g564(.A(new_n239), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT107), .B1(new_n663), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n687), .A2(new_n748), .A3(new_n702), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n590), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n731), .A2(new_n755), .A3(new_n733), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  AOI211_X1 g572(.A(new_n667), .B(new_n744), .C1(new_n746), .C2(new_n747), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n740), .A2(new_n759), .A3(new_n717), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NAND2_X1  g575(.A1(new_n441), .A2(new_n377), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n437), .B2(new_n439), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT108), .B1(new_n479), .B2(new_n481), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n609), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n766), .A3(G469), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n487), .A3(new_n612), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n763), .A2(new_n605), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n372), .A2(new_n374), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n698), .A2(KEYINPUT32), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n753), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n629), .A2(KEYINPUT42), .A3(new_n641), .A4(new_n679), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n774), .A3(KEYINPUT109), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n347), .B1(new_n343), .B2(new_n345), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n372), .A3(new_n374), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n753), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n763), .A2(new_n605), .A3(new_n768), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT42), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n357), .B1(new_n725), .B2(new_n726), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n449), .B1(new_n784), .B2(new_n448), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n447), .B1(new_n785), .B2(new_n767), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n683), .A2(new_n786), .A3(new_n606), .A4(new_n763), .ZN(new_n787));
  INV_X1    g601(.A(new_n717), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT110), .B(G131), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G33));
  NAND2_X1  g606(.A1(new_n680), .A2(new_n681), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n769), .A2(new_n795), .A3(new_n376), .A4(new_n682), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  XNOR2_X1  g612(.A(new_n701), .B(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n641), .A2(KEYINPUT43), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n629), .A2(new_n640), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n799), .A2(new_n800), .B1(KEYINPUT43), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n617), .A2(new_n667), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT113), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n802), .A2(new_n807), .A3(KEYINPUT44), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n482), .A2(KEYINPUT45), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n448), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n764), .A2(new_n766), .A3(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n449), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT46), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n487), .B1(new_n813), .B2(KEYINPUT46), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n605), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n763), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n804), .B2(new_n805), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n706), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n816), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n788), .A2(new_n683), .A3(new_n606), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n763), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  NAND3_X1  g640(.A1(new_n641), .A2(new_n377), .A3(new_n605), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n827), .B(new_n799), .C1(new_n752), .C2(new_n750), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n723), .A2(new_n729), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT49), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n692), .A3(new_n700), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n748), .A2(new_n753), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n802), .A2(new_n676), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n730), .A2(new_n377), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n692), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n692), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n833), .A2(new_n836), .A3(KEYINPUT50), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n829), .A2(new_n447), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n763), .B(new_n833), .C1(new_n823), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n818), .A2(new_n730), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n240), .A2(new_n674), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n700), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n629), .A3(new_n641), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n802), .A2(new_n676), .A3(new_n846), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n759), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(KEYINPUT115), .A3(new_n853), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT51), .A4(new_n851), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n740), .ZN(new_n859));
  INV_X1    g673(.A(new_n645), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n859), .B(new_n589), .C1(new_n860), .C2(new_n848), .ZN(new_n861));
  INV_X1    g675(.A(new_n772), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT48), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(KEYINPUT48), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n782), .A2(new_n789), .B1(new_n794), .B2(new_n796), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n741), .A2(new_n592), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n423), .A2(new_n438), .A3(new_n435), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n438), .B1(new_n423), .B2(new_n435), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n379), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n377), .B1(new_n873), .B2(new_n626), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n629), .A2(new_n640), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n755), .A3(new_n584), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n621), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n376), .A2(new_n731), .A3(new_n733), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n628), .A2(new_n582), .A3(new_n672), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n748), .A2(new_n702), .A3(new_n687), .A4(new_n753), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n731), .A2(new_n755), .A3(new_n733), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n879), .A2(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n628), .B1(new_n642), .B2(new_n644), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n669), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n759), .A2(new_n717), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n685), .B1(new_n356), .B2(new_n375), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n583), .A2(new_n763), .A3(new_n672), .A4(new_n679), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n887), .A2(new_n769), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n869), .A2(new_n878), .A3(new_n886), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n667), .A2(new_n679), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n356), .B2(new_n699), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n687), .A3(new_n702), .A4(new_n786), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n688), .A2(new_n760), .A3(new_n718), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n888), .B(new_n687), .C1(new_n682), .C2(new_n717), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT52), .A3(new_n760), .A4(new_n894), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n868), .B1(new_n891), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n735), .A2(new_n757), .A3(new_n738), .A4(new_n669), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n615), .A2(new_n620), .A3(new_n877), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n592), .A3(new_n741), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n769), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n889), .A2(new_n888), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n902), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n897), .A2(new_n899), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(KEYINPUT53), .A3(new_n909), .A4(new_n869), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n901), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n901), .A2(new_n910), .A3(KEYINPUT54), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n867), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(G952), .A2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n831), .B1(new_n915), .B2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n221), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n226), .B1(new_n901), .B2(new_n910), .ZN(new_n920));
  INV_X1    g734(.A(new_n379), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n410), .B1(new_n419), .B2(new_n422), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n415), .ZN(new_n924));
  XOR2_X1   g738(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n920), .A2(KEYINPUT117), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n920), .A2(KEYINPUT117), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n921), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n931), .B2(new_n933), .ZN(G51));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n812), .A3(new_n811), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n449), .B(KEYINPUT57), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n913), .A2(new_n914), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n727), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n918), .B1(new_n935), .B2(new_n938), .ZN(G54));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n536), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n928), .A2(new_n929), .A3(new_n652), .A4(new_n940), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n918), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n913), .A2(new_n914), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n634), .A2(new_n637), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT118), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n947), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n919), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n913), .A2(new_n914), .A3(new_n950), .A4(new_n946), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT123), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n911), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(KEYINPUT121), .A3(new_n665), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n919), .B1(new_n959), .B2(KEYINPUT61), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n965), .B2(new_n236), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT121), .B1(new_n966), .B2(new_n665), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n961), .A3(new_n967), .A4(new_n969), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n588), .B2(new_n413), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n902), .A2(new_n904), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n923), .B1(G898), .B2(new_n221), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  AOI21_X1  g794(.A(new_n221), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n365), .A2(new_n337), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n529), .A2(new_n530), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n862), .A2(new_n687), .A3(new_n702), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n817), .A2(new_n706), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n898), .A2(new_n760), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n869), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n820), .A2(new_n825), .A3(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n984), .B(new_n985), .C1(new_n990), .C2(G953), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n875), .A2(new_n584), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n708), .A2(new_n376), .A3(new_n763), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n820), .A2(new_n825), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT103), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n714), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n714), .A2(new_n996), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n998), .A3(new_n988), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n715), .A2(new_n1001), .A3(new_n988), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n984), .B1(new_n1003), .B2(new_n221), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n981), .B1(new_n992), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n991), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n981), .B(KEYINPUT124), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(G72));
  XOR2_X1   g823(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1010));
  NOR2_X1   g824(.A1(new_n598), .A2(new_n446), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n977), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1003), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n694), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1012), .B1(new_n990), .B2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n368), .A2(new_n246), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n918), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n694), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT127), .B1(new_n911), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n911), .A2(KEYINPUT127), .A3(new_n1021), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1016), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(G57));
endmodule


