

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XNOR2_X1 U324 ( .A(n415), .B(n350), .ZN(n351) );
  XOR2_X1 U325 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XNOR2_X1 U326 ( .A(n352), .B(n351), .ZN(n354) );
  NAND2_X1 U327 ( .A1(n567), .A2(n459), .ZN(n426) );
  XNOR2_X1 U328 ( .A(n426), .B(KEYINPUT55), .ZN(n443) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n444) );
  XOR2_X1 U330 ( .A(n358), .B(n357), .Z(n541) );
  XNOR2_X1 U331 ( .A(n444), .B(KEYINPUT58), .ZN(n445) );
  XNOR2_X1 U332 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  XNOR2_X1 U333 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n292), .B(n293), .ZN(n352) );
  XNOR2_X1 U335 ( .A(G50GAT), .B(KEYINPUT71), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n294), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U337 ( .A(n352), .B(n409), .ZN(n307) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G85GAT), .Z(n360) );
  XOR2_X1 U339 ( .A(G36GAT), .B(G190GAT), .Z(n400) );
  XOR2_X1 U340 ( .A(n360), .B(n400), .Z(n296) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U343 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n298) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(G92GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT74), .Z(n309) );
  XOR2_X1 U348 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n302) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n309), .B(n303), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n307), .B(n306), .Z(n464) );
  XNOR2_X1 U354 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n308), .B(KEYINPUT3), .ZN(n420) );
  XOR2_X1 U356 ( .A(n309), .B(n420), .Z(n311) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(n312), .B(KEYINPUT87), .Z(n315) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n313), .B(G120GAT), .ZN(n438) );
  XNOR2_X1 U362 ( .A(n438), .B(KEYINPUT5), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G162GAT), .Z(n317) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(G127GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U367 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n321) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT86), .B(KEYINPUT6), .Z(n323) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U375 ( .A(n327), .B(n326), .Z(n457) );
  XNOR2_X1 U376 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n388) );
  INV_X1 U377 ( .A(n464), .ZN(n551) );
  XOR2_X1 U378 ( .A(KEYINPUT76), .B(G64GAT), .Z(n329) );
  XNOR2_X1 U379 ( .A(G22GAT), .B(G78GAT), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n343) );
  XOR2_X1 U385 ( .A(G1GAT), .B(KEYINPUT64), .Z(n353) );
  XNOR2_X1 U386 ( .A(G71GAT), .B(G57GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(KEYINPUT13), .ZN(n359) );
  XOR2_X1 U388 ( .A(n359), .B(KEYINPUT75), .Z(n336) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n353), .B(n337), .ZN(n341) );
  XOR2_X1 U392 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XOR2_X1 U393 ( .A(n396), .B(G155GAT), .Z(n339) );
  XOR2_X1 U394 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XNOR2_X1 U395 ( .A(n434), .B(G211GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U398 ( .A(n343), .B(n342), .Z(n576) );
  INV_X1 U399 ( .A(n576), .ZN(n548) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G113GAT), .Z(n345) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U403 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n347) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n358) );
  XOR2_X1 U407 ( .A(G141GAT), .B(G22GAT), .Z(n415) );
  AND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n356) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U412 ( .A(n541), .ZN(n568) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(n359), .Z(n362) );
  XNOR2_X1 U414 ( .A(G120GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n367) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n363), .B(G148GAT), .ZN(n418) );
  XOR2_X1 U418 ( .A(n418), .B(KEYINPUT32), .Z(n365) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U421 ( .A(n367), .B(n366), .Z(n375) );
  XOR2_X1 U422 ( .A(G92GAT), .B(KEYINPUT68), .Z(n369) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(G64GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(G204GAT), .B(n370), .Z(n395) );
  XOR2_X1 U426 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT33), .B(KEYINPUT66), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n395), .B(n373), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n573) );
  XNOR2_X1 U431 ( .A(n573), .B(KEYINPUT41), .ZN(n543) );
  INV_X1 U432 ( .A(n543), .ZN(n557) );
  NOR2_X1 U433 ( .A1(n568), .A2(n557), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n376), .B(KEYINPUT46), .ZN(n377) );
  NOR2_X1 U435 ( .A1(n548), .A2(n377), .ZN(n378) );
  XOR2_X1 U436 ( .A(n378), .B(KEYINPUT110), .Z(n379) );
  NOR2_X2 U437 ( .A1(n551), .A2(n379), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n380), .B(KEYINPUT47), .ZN(n386) );
  XNOR2_X1 U439 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n381) );
  XOR2_X1 U440 ( .A(n381), .B(n551), .Z(n579) );
  NOR2_X1 U441 ( .A1(n579), .A2(n576), .ZN(n382) );
  XOR2_X1 U442 ( .A(KEYINPUT45), .B(n382), .Z(n383) );
  NOR2_X1 U443 ( .A1(n541), .A2(n383), .ZN(n384) );
  NAND2_X1 U444 ( .A1(n384), .A2(n573), .ZN(n385) );
  NAND2_X1 U445 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n540) );
  XOR2_X1 U447 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n390) );
  XNOR2_X1 U448 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U450 ( .A(G169GAT), .B(n391), .Z(n430) );
  XOR2_X1 U451 ( .A(KEYINPUT83), .B(G218GAT), .Z(n393) );
  XNOR2_X1 U452 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U454 ( .A(G197GAT), .B(n394), .Z(n421) );
  XNOR2_X1 U455 ( .A(n421), .B(n395), .ZN(n404) );
  XOR2_X1 U456 ( .A(n396), .B(KEYINPUT90), .Z(n398) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U459 ( .A(n399), .B(KEYINPUT88), .Z(n402) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT89), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(n430), .B(n405), .Z(n511) );
  INV_X1 U464 ( .A(n511), .ZN(n406) );
  NOR2_X1 U465 ( .A1(n540), .A2(n406), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n407), .B(KEYINPUT54), .ZN(n408) );
  AND2_X1 U467 ( .A1(n457), .A2(n408), .ZN(n567) );
  XOR2_X1 U468 ( .A(n409), .B(KEYINPUT22), .Z(n411) );
  NAND2_X1 U469 ( .A1(G228GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n425) );
  XOR2_X1 U471 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U472 ( .A(G204GAT), .B(KEYINPUT85), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U474 ( .A(n414), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U475 ( .A(n415), .B(KEYINPUT84), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n459) );
  XOR2_X1 U481 ( .A(KEYINPUT79), .B(G176GAT), .Z(n428) );
  XNOR2_X1 U482 ( .A(KEYINPUT80), .B(G71GAT), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U485 ( .A(G134GAT), .B(G190GAT), .Z(n432) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G99GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n437), .B(G183GAT), .Z(n440) );
  XNOR2_X1 U492 ( .A(n438), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n522) );
  NAND2_X1 U495 ( .A1(n443), .A2(n522), .ZN(n563) );
  NOR2_X1 U496 ( .A1(n464), .A2(n563), .ZN(n446) );
  NAND2_X1 U497 ( .A1(n541), .A2(n573), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(KEYINPUT70), .ZN(n485) );
  NAND2_X1 U499 ( .A1(n511), .A2(n522), .ZN(n448) );
  NAND2_X1 U500 ( .A1(n448), .A2(n459), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n449), .B(KEYINPUT25), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT94), .B(n450), .Z(n455) );
  XNOR2_X1 U503 ( .A(KEYINPUT93), .B(KEYINPUT26), .ZN(n452) );
  NOR2_X1 U504 ( .A1(n522), .A2(n459), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U506 ( .A(KEYINPUT92), .B(n453), .Z(n566) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(n511), .ZN(n458) );
  NAND2_X1 U508 ( .A1(n566), .A2(n458), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n456), .A2(n457), .ZN(n463) );
  INV_X1 U511 ( .A(n457), .ZN(n509) );
  AND2_X1 U512 ( .A1(n458), .A2(n509), .ZN(n538) );
  XOR2_X1 U513 ( .A(n459), .B(KEYINPUT28), .Z(n517) );
  INV_X1 U514 ( .A(n517), .ZN(n460) );
  NAND2_X1 U515 ( .A1(n538), .A2(n460), .ZN(n521) );
  NOR2_X1 U516 ( .A1(n522), .A2(n521), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT91), .B(n461), .ZN(n462) );
  NAND2_X1 U518 ( .A1(n463), .A2(n462), .ZN(n480) );
  XOR2_X1 U519 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n466) );
  NAND2_X1 U520 ( .A1(n548), .A2(n464), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n480), .A2(n467), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT95), .B(n468), .Z(n496) );
  NOR2_X1 U524 ( .A1(n485), .A2(n496), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT96), .B(n469), .ZN(n478) );
  NAND2_X1 U526 ( .A1(n478), .A2(n509), .ZN(n473) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n471) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n473), .B(n472), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT99), .Z(n475) );
  NAND2_X1 U532 ( .A1(n511), .A2(n478), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U535 ( .A1(n522), .A2(n478), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NAND2_X1 U537 ( .A1(n478), .A2(n517), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n489) );
  INV_X1 U540 ( .A(KEYINPUT101), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n576), .A2(n480), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n579), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n484), .ZN(n506) );
  NOR2_X1 U545 ( .A1(n485), .A2(n506), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n494) );
  NAND2_X1 U548 ( .A1(n494), .A2(n509), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U550 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U551 ( .A1(n494), .A2(n511), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n494), .A2(n522), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n494), .A2(n517), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n499) );
  NAND2_X1 U559 ( .A1(n568), .A2(n543), .ZN(n507) );
  NOR2_X1 U560 ( .A1(n507), .A2(n496), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(n497), .Z(n503) );
  NAND2_X1 U562 ( .A1(n503), .A2(n509), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n511), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n503), .A2(n522), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U570 ( .A1(n503), .A2(n517), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(KEYINPUT106), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n509), .A2(n516), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  XOR2_X1 U576 ( .A(G92GAT), .B(KEYINPUT107), .Z(n513) );
  NAND2_X1 U577 ( .A1(n511), .A2(n516), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n522), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G99GAT), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n526) );
  NOR2_X1 U587 ( .A1(n540), .A2(n521), .ZN(n523) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(n524), .Z(n534) );
  NAND2_X1 U590 ( .A1(n534), .A2(n541), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U594 ( .A1(n534), .A2(n543), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT115), .Z(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n548), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n551), .A2(n534), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n537), .Z(G1343GAT) );
  NAND2_X1 U605 ( .A1(n566), .A2(n538), .ZN(n539) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n541), .A2(n552), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n545) );
  NAND2_X1 U611 ( .A1(n552), .A2(n543), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U615 ( .A1(n552), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n568), .A2(n563), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT56), .B(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U629 ( .A1(n576), .A2(n563), .ZN(n564) );
  XOR2_X1 U630 ( .A(n564), .B(KEYINPUT124), .Z(n565) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n578), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n578), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(G218GAT), .B(n582), .Z(G1355GAT) );
endmodule

