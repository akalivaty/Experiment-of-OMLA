//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(KEYINPUT67), .B1(G567), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n466), .B2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n467), .C2(new_n466), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(G2104), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n497), .B1(new_n496), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(G164));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT71), .B(G88), .Z(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g093(.A(G50), .B(G543), .C1(new_n508), .C2(new_n507), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n514), .A2(KEYINPUT69), .A3(G50), .A4(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n509), .A2(new_n510), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n523), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND3_X1   g105(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT7), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n514), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI211_X1 g110(.A(new_n531), .B(new_n533), .C1(G51), .C2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n512), .A2(new_n516), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G651), .B1(G52), .B2(new_n535), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n512), .A2(new_n516), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n537), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(G43), .A2(new_n535), .B1(new_n550), .B2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n535), .A2(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(KEYINPUT73), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n561), .B(KEYINPUT9), .C1(new_n559), .C2(new_n560), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n559), .B(new_n563), .C1(new_n560), .C2(KEYINPUT73), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G651), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n537), .A2(G91), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n562), .A2(new_n564), .A3(new_n567), .A4(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n566), .B1(new_n525), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n535), .B2(G49), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n544), .ZN(G288));
  OAI21_X1  g150(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n513), .A2(KEYINPUT74), .A3(G61), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n512), .A2(G86), .A3(new_n516), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n535), .A2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n535), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n566), .B2(new_n588), .C1(new_n544), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT75), .Z(new_n592));
  NAND2_X1  g167(.A1(new_n537), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n525), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(G54), .A2(new_n535), .B1(new_n598), .B2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AND4_X1   g179(.A1(new_n562), .A2(new_n564), .A3(new_n567), .A4(new_n568), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XNOR2_X1  g182(.A(KEYINPUT76), .B(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(G860), .B2(new_n608), .ZN(G148));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n553), .ZN(G323));
  XOR2_X1   g187(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  NAND2_X1  g189(.A1(new_n477), .A2(new_n473), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n484), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n465), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n479), .A2(KEYINPUT78), .A3(G123), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n479), .B2(G123), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n619), .B1(new_n620), .B2(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n618), .A2(G2100), .B1(G2096), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n625), .B(new_n627), .C1(G2096), .C2(new_n624), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT79), .Z(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n626), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n647), .A2(new_n648), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  OR2_X1    g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n665), .A3(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n665), .C2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT33), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1976), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(G16), .A2(G22), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G166), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT85), .B(G1971), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT83), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n484), .A2(G131), .ZN(new_n697));
  INV_X1    g272(.A(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n478), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n693), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT84), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n704), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n691), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT86), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT86), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n682), .A2(new_n686), .A3(new_n690), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n713), .A2(new_n714), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n711), .B2(new_n712), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n718), .B1(new_n721), .B2(KEYINPUT88), .ZN(new_n722));
  NAND2_X1  g297(.A1(G168), .A2(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(KEYINPUT93), .C1(G16), .C2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT93), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1966), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2072), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT25), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G139), .B2(new_n484), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT90), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n465), .B2(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G33), .B(new_n735), .S(G29), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n728), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n729), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n677), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT23), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n605), .B2(new_n677), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n677), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n601), .B2(new_n677), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n692), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n692), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(G1348), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n747), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2090), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n692), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n484), .A2(G140), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT89), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(G116), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n479), .B2(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n758), .B(new_n769), .C1(G1966), .C2(new_n725), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n473), .A2(G105), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n479), .A2(G129), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n484), .A2(G141), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  AND4_X1   g350(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(new_n692), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n692), .B2(G32), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(G34), .ZN(new_n782));
  INV_X1    g357(.A(G160), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(G2084), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g362(.A1(G5), .A2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT96), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G301), .B2(new_n677), .ZN(new_n790));
  INV_X1    g365(.A(G1961), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT95), .B(G28), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(new_n692), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n793), .B1(new_n795), .B2(new_n797), .C1(new_n624), .C2(new_n692), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n778), .B2(new_n779), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n786), .A2(new_n787), .A3(new_n792), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n553), .A2(new_n677), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n677), .B2(G19), .ZN(new_n802));
  INV_X1    g377(.A(G1341), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n790), .A2(new_n791), .ZN(new_n805));
  INV_X1    g380(.A(new_n802), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G1341), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n770), .A2(new_n800), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n738), .A2(new_n744), .A3(new_n753), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n721), .B2(new_n717), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n720), .A2(new_n722), .A3(new_n810), .ZN(G311));
  NAND3_X1  g386(.A1(new_n720), .A2(new_n722), .A3(new_n810), .ZN(G150));
  AND3_X1   g387(.A1(new_n512), .A2(G93), .A3(new_n516), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n814), .A2(new_n566), .B1(new_n815), .B2(new_n534), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT37), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n601), .A2(G559), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n552), .A2(new_n817), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT101), .ZN(new_n826));
  INV_X1    g401(.A(new_n817), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n553), .A2(new_n827), .A3(KEYINPUT100), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n552), .B2(new_n817), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n824), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n836), .A3(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n821), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g417(.A(KEYINPUT102), .B(KEYINPUT39), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n818), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n820), .B1(new_n844), .B2(new_n845), .ZN(G145));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n496), .A2(new_n503), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n767), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n735), .ZN(new_n850));
  INV_X1    g425(.A(new_n776), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n700), .B(new_n616), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n484), .A2(G142), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n465), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  INV_X1    g431(.A(G130), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n854), .B1(new_n855), .B2(new_n856), .C1(new_n857), .C2(new_n478), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n853), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n488), .B(new_n783), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n624), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n859), .B(KEYINPUT103), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n860), .B(new_n863), .C1(new_n852), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n852), .Z(new_n866));
  OAI211_X1 g441(.A(new_n847), .B(new_n865), .C1(new_n866), .C2(new_n863), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g443(.A1(new_n605), .A2(new_n595), .A3(new_n599), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n600), .A2(G299), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n832), .B(new_n610), .ZN(new_n878));
  MUX2_X1   g453(.A(new_n871), .B(new_n877), .S(new_n878), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n679), .B(G305), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(G166), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n880), .B(new_n881), .Z(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT42), .Z(new_n883));
  XOR2_X1   g458(.A(new_n879), .B(new_n883), .Z(new_n884));
  MUX2_X1   g459(.A(new_n827), .B(new_n884), .S(G868), .Z(G295));
  MUX2_X1   g460(.A(new_n827), .B(new_n884), .S(G868), .Z(G331));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n826), .A2(new_n831), .A3(G301), .ZN(new_n888));
  AOI21_X1  g463(.A(G301), .B1(new_n826), .B2(new_n831), .ZN(new_n889));
  OAI21_X1  g464(.A(G286), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n832), .A2(G171), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n826), .A2(new_n831), .A3(G301), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(G168), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n893), .A3(new_n871), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n869), .B2(new_n870), .ZN(new_n897));
  INV_X1    g472(.A(new_n874), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n871), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n894), .A2(new_n895), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n890), .A2(new_n893), .A3(new_n871), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n887), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n896), .A2(new_n877), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n887), .A3(new_n894), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n847), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n876), .B1(new_n890), .B2(new_n893), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n887), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n882), .B1(new_n901), .B2(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT43), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n903), .A2(new_n906), .A3(KEYINPUT43), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n918), .ZN(G397));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(G160), .B2(G40), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n484), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n922));
  INV_X1    g497(.A(G125), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n482), .B2(new_n483), .ZN(new_n924));
  INV_X1    g499(.A(new_n469), .ZN(new_n925));
  OAI21_X1  g500(.A(G2105), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND4_X1   g501(.A1(KEYINPUT107), .A2(new_n922), .A3(new_n926), .A4(G40), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n848), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n920), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n922), .A2(new_n926), .A3(G40), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(G160), .A2(KEYINPUT107), .A3(G40), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n938), .A2(KEYINPUT108), .A3(new_n930), .A4(new_n931), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT109), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n776), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(G1996), .A3(new_n851), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(KEYINPUT110), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n767), .B(G2067), .Z(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n946), .A2(new_n947), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n696), .A2(new_n704), .A3(new_n699), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n700), .A2(new_n703), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n940), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  AND2_X1   g529(.A1(G290), .A2(G1986), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n940), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n944), .A2(new_n950), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT111), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT116), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n848), .B2(new_n929), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT112), .B(G1384), .C1(new_n496), .C2(new_n503), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n959), .B(new_n938), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n921), .B2(new_n927), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n498), .A2(new_n502), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n493), .B2(new_n495), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n968), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(new_n495), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n494), .B1(new_n477), .B2(new_n491), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n960), .B(new_n929), .C1(new_n972), .C2(new_n967), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT116), .B(new_n966), .C1(new_n974), .C2(new_n928), .ZN(new_n975));
  INV_X1    g550(.A(G2090), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n848), .A2(KEYINPUT68), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n497), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n964), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n965), .A2(new_n975), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n929), .B1(new_n504), .B2(new_n505), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n931), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n968), .A2(G1384), .ZN(new_n984));
  AOI22_X1  g559(.A1(KEYINPUT45), .A2(new_n984), .B1(new_n936), .B2(new_n937), .ZN(new_n985));
  AOI21_X1  g560(.A(G1971), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G8), .ZN(new_n989));
  NAND3_X1  g564(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n991), .B2(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(new_n992), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(KEYINPUT114), .A3(new_n990), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n938), .A2(new_n976), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n969), .A2(new_n964), .A3(new_n973), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(KEYINPUT113), .C1(new_n979), .C2(new_n964), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n982), .A2(new_n1003), .A3(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n999), .B(G8), .C1(new_n1005), .C2(new_n986), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n938), .A2(new_n969), .A3(new_n973), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n679), .A2(G1976), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(G8), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1007), .A2(G8), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n584), .A2(new_n585), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n576), .A2(new_n577), .B1(G73), .B2(G543), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n566), .B1(new_n1016), .B2(new_n581), .ZN(new_n1017));
  OAI21_X1  g592(.A(G1981), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n583), .A2(new_n1019), .A3(new_n584), .A4(new_n585), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1020), .A3(KEYINPUT49), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1007), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT115), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1007), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1024), .A4(new_n1023), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1014), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n994), .A2(KEYINPUT125), .A3(new_n1006), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT125), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1014), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1006), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n993), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n988), .B2(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1966), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n931), .A2(G1384), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n938), .B1(G164), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n969), .B2(new_n973), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT117), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n928), .A2(G2084), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G168), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1046), .A3(G168), .A4(new_n1047), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(new_n938), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT122), .B(G1961), .Z(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n928), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1062), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(KEYINPUT123), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G2078), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n922), .A2(G40), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n924), .A2(new_n925), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n465), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n932), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n983), .A2(new_n750), .A3(new_n985), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1079), .B2(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(G171), .B1(new_n1067), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1082), .A2(new_n1069), .B1(new_n1078), .B2(new_n1068), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(G301), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(KEYINPUT126), .A3(G301), .A4(new_n1083), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(new_n1089), .A3(KEYINPUT54), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1061), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT123), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1093));
  AOI211_X1 g668(.A(G171), .B(new_n1080), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G301), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1039), .A2(new_n1059), .A3(new_n1090), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n605), .B(KEYINPUT57), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n965), .A2(new_n975), .A3(new_n980), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n983), .A2(new_n985), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1099), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT120), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1099), .B(new_n1108), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1098), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1099), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1098), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1104), .A2(new_n1118), .A3(new_n1099), .A4(new_n1108), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1112), .A2(KEYINPUT121), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1007), .A2(G2067), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1061), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n601), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1106), .A2(new_n941), .ZN(new_n1128));
  OR2_X1    g703(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1129));
  NAND2_X1  g704(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1007), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1132), .B2(new_n553), .ZN(new_n1133));
  AOI211_X1 g708(.A(KEYINPUT59), .B(new_n552), .C1(new_n1128), .C2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1126), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1124), .B(new_n600), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(KEYINPUT60), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1114), .A2(new_n1121), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1124), .A2(new_n600), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1112), .B1(new_n1109), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1097), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1031), .A2(new_n1038), .A3(new_n1095), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1051), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1144));
  OAI21_X1  g719(.A(G286), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1057), .B1(new_n1056), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1054), .A2(KEYINPUT51), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT62), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1055), .A2(new_n1149), .A3(new_n1058), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1142), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1006), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  NAND2_X1  g728(.A1(G168), .A2(G8), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .A4(new_n994), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1159), .B2(new_n1155), .ZN(new_n1160));
  OAI21_X1  g735(.A(G8), .B1(new_n1005), .B2(new_n986), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n993), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1162), .A2(new_n1030), .A3(KEYINPUT119), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1030), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1155), .A2(KEYINPUT63), .A3(new_n1006), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1158), .A2(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1033), .A2(new_n1011), .A3(new_n679), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1020), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1006), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1169), .A2(new_n1027), .B1(new_n1170), .B2(new_n1030), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1151), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n958), .B1(new_n1141), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n940), .B1(new_n949), .B2(new_n851), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT46), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n943), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n943), .A2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT47), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT47), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1180), .B(new_n1174), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n944), .A2(new_n950), .A3(new_n953), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n944), .A2(KEYINPUT127), .A3(new_n950), .A4(new_n953), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n940), .A2(new_n954), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT48), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n767), .A2(G2067), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n940), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1182), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1173), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g769(.A1(G227), .A2(new_n463), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1196), .A2(new_n644), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G229), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g772(.A(new_n867), .B(new_n1198), .C1(new_n916), .C2(new_n917), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


