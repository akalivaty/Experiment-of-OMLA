//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n205), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n219), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n250), .A2(new_n215), .A3(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n214), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G50), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n250), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(G50), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT8), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n268), .B1(G150), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n203), .A2(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n261), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n260), .B1(KEYINPUT69), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(KEYINPUT69), .B2(new_n272), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n274), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT72), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n267), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(KEYINPUT68), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  INV_X1    g0090(.A(new_n287), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(G1698), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n289), .B1(new_n290), .B2(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  OAI211_X1 g0097(.A(G1), .B(G13), .C1(new_n267), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G274), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n295), .A2(new_n300), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT67), .B(G226), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(G200), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n278), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT73), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n311), .A2(G190), .B1(new_n275), .B2(new_n274), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n309), .A2(new_n310), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n314), .A2(new_n313), .A3(new_n278), .A4(new_n308), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n274), .C1(G179), .C2(new_n306), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n282), .A2(new_n286), .A3(G226), .A4(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n282), .A2(new_n286), .A3(G232), .A4(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n295), .ZN(new_n328));
  INV_X1    g0128(.A(new_n300), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n298), .ZN(new_n330));
  INV_X1    g0130(.A(G238), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n301), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n327), .B2(new_n295), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT74), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(G169), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(new_n343), .A3(G169), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n337), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n335), .A2(G179), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n254), .A2(G68), .A3(new_n256), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT12), .ZN(new_n349));
  INV_X1    g0149(.A(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n251), .B2(new_n350), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n354), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n268), .A2(G77), .B1(G20), .B2(new_n350), .ZN(new_n357));
  NOR4_X1   g0157(.A1(new_n202), .A2(KEYINPUT75), .A3(G20), .A4(G33), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n269), .B2(G50), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n357), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n361), .A2(new_n362), .A3(new_n253), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n361), .B2(new_n253), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n355), .A2(new_n356), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n347), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n339), .A2(G200), .A3(new_n340), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n334), .B2(KEYINPUT13), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n365), .B1(new_n345), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n254), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n266), .A2(new_n256), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(new_n259), .B2(new_n266), .ZN(new_n376));
  AND2_X1   g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT77), .B(G20), .C1(new_n377), .C2(new_n201), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n269), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(G58), .B(G68), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT77), .B1(new_n381), .B2(G20), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT78), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n280), .A2(new_n281), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(new_n215), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n280), .A2(new_n281), .A3(new_n386), .A4(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n377), .B2(new_n201), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT78), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n379), .A4(new_n378), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n383), .A2(new_n388), .A3(KEYINPUT16), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n253), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n280), .A2(new_n281), .A3(new_n279), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT68), .B1(new_n284), .B2(new_n285), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n215), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n386), .ZN(new_n400));
  INV_X1    g0200(.A(new_n387), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n350), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n383), .A2(new_n393), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n395), .B1(new_n404), .B2(KEYINPUT79), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n383), .A2(new_n393), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n282), .B2(new_n286), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n401), .B1(new_n407), .B2(KEYINPUT7), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G68), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT16), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT79), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n376), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n303), .A2(G232), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n301), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n284), .A2(new_n285), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n292), .A2(new_n323), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(G226), .C2(new_n323), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n298), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(new_n414), .A3(new_n301), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G179), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n423), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n425), .A2(new_n421), .A3(new_n416), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n319), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n413), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n376), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n394), .A2(new_n253), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n410), .B2(new_n411), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n404), .A2(KEYINPUT79), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n427), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n422), .A2(new_n368), .A3(new_n423), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n426), .B2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n430), .B(new_n440), .C1(new_n432), .C2(new_n433), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G244), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n301), .B1(new_n330), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n288), .A2(G232), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n450), .B1(new_n206), .B2(new_n291), .C1(new_n293), .C2(new_n331), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(new_n295), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n266), .B1(KEYINPUT70), .B2(new_n269), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(KEYINPUT70), .B2(new_n269), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  INV_X1    g0255(.A(new_n268), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n455), .A2(new_n456), .B1(new_n215), .B2(new_n290), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n253), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT71), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n254), .A2(G77), .A3(new_n256), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G77), .B2(new_n259), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n452), .A2(G169), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G179), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n459), .A2(new_n461), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n452), .A2(G190), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n468), .C1(new_n312), .C2(new_n452), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR4_X1   g0270(.A1(new_n322), .A2(new_n373), .A3(new_n447), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n331), .A2(new_n323), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n448), .A2(G1698), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n280), .C2(new_n281), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT84), .A2(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT84), .A2(G116), .ZN(new_n476));
  OAI21_X1  g0276(.A(G33), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n298), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n299), .A2(G1), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n222), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n298), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n298), .A2(G274), .ZN(new_n486));
  INV_X1    g0286(.A(new_n483), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT86), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n474), .A2(new_n480), .A3(new_n477), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n474), .B2(new_n477), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n295), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n488), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n463), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT19), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n456), .B2(new_n205), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n417), .A2(new_n215), .A3(G68), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n215), .B1(new_n326), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(G87), .B2(new_n207), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n253), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n455), .A2(new_n251), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n255), .A2(KEYINPUT83), .A3(G33), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n267), .B2(G1), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n261), .A2(new_n259), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n503), .B(new_n504), .C1(new_n455), .C2(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n488), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n494), .B1(new_n492), .B2(new_n493), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n496), .B(new_n509), .C1(new_n512), .C2(G169), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n489), .A2(G190), .A3(new_n495), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n503), .A2(new_n504), .ZN(new_n515));
  INV_X1    g0315(.A(new_n508), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(G87), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n514), .B(new_n517), .C1(new_n512), .C2(new_n312), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n298), .A3(G274), .A4(new_n483), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n483), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n298), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n520), .B1(new_n524), .B2(new_n223), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n282), .A2(new_n286), .A3(G250), .A4(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n448), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n282), .A2(new_n286), .A3(new_n323), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(new_n323), .C1(new_n280), .C2(new_n281), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n527), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n526), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n525), .B1(new_n533), .B2(new_n295), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n319), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n259), .B2(G97), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n205), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n516), .A2(G97), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  NOR2_X1   g0341(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n542), .B1(KEYINPUT6), .B2(new_n205), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(G20), .C1(new_n541), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n269), .A2(G77), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(G107), .B2(new_n408), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n540), .B1(new_n549), .B2(new_n261), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n534), .A2(new_n463), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n536), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n534), .A2(new_n368), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G200), .B2(new_n534), .ZN(new_n554));
  INV_X1    g0354(.A(new_n540), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n408), .A2(G107), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n547), .A3(new_n546), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n557), .B2(new_n253), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n513), .A2(new_n518), .A3(new_n552), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n223), .A2(new_n323), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n417), .A2(new_n561), .B1(G33), .B2(G294), .ZN(new_n562));
  OAI211_X1 g0362(.A(G250), .B(new_n323), .C1(new_n280), .C2(new_n281), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n417), .A2(new_n565), .A3(G250), .A4(new_n323), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n295), .ZN(new_n568));
  INV_X1    g0368(.A(new_n524), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G264), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n520), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT90), .B1(new_n571), .B2(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n312), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n567), .A2(new_n295), .B1(G264), .B2(new_n569), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT90), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n368), .A4(new_n520), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n417), .A2(new_n215), .A3(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n221), .A2(KEYINPUT22), .A3(G20), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n282), .A2(new_n286), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n477), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n215), .B2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n583), .A2(new_n215), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT24), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n261), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n259), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n516), .A2(G107), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n577), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n574), .A2(new_n463), .A3(new_n520), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n571), .A2(new_n319), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n592), .C2(new_n597), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n475), .A2(new_n476), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G20), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n605), .A2(G1), .A3(new_n250), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n530), .B(new_n215), .C1(G33), .C2(new_n205), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT84), .B(G116), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n253), .B(new_n607), .C1(new_n608), .C2(new_n215), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n605), .A2(KEYINPUT20), .A3(new_n607), .A4(new_n253), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT88), .B1(new_n508), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n507), .A2(new_n505), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n254), .A2(new_n616), .A3(new_n617), .A4(G116), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n223), .A2(new_n323), .ZN(new_n621));
  OAI221_X1 g0421(.A(new_n621), .B1(G264), .B2(new_n323), .C1(new_n280), .C2(new_n281), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G303), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n282), .B2(new_n286), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n295), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n523), .A2(G270), .A3(new_n298), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n627), .A2(new_n520), .A3(KEYINPUT87), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT87), .B1(new_n627), .B2(new_n520), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n620), .A2(G169), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n613), .A2(new_n619), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n626), .B(G179), .C1(new_n628), .C2(new_n629), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(G200), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n634), .C1(new_n368), .C2(new_n630), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n620), .A2(KEYINPUT21), .A3(G169), .A4(new_n630), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n633), .A2(new_n636), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n560), .A2(new_n603), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n471), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n642), .B(KEYINPUT91), .Z(G372));
  NOR2_X1   g0443(.A1(new_n482), .A2(new_n488), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n496), .B(new_n509), .C1(G169), .C2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n514), .B(new_n517), .C1(new_n312), .C2(new_n644), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n599), .A2(new_n552), .A3(new_n559), .A4(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n636), .A2(new_n639), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n602), .A3(new_n633), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n536), .A2(new_n550), .A3(new_n551), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n647), .A3(new_n645), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n513), .A2(new_n518), .A3(new_n652), .A4(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n471), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n372), .A2(new_n465), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n445), .B1(new_n660), .B2(new_n366), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n318), .B1(new_n661), .B2(new_n437), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n321), .A3(new_n662), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n649), .A2(new_n633), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n258), .A2(new_n215), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n634), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n640), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n591), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n590), .B1(new_n582), .B2(new_n587), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n253), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(new_n596), .B1(new_n319), .B2(new_n571), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(new_n600), .B1(new_n577), .B2(new_n598), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n598), .B2(new_n671), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n602), .B2(new_n671), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n682), .A2(new_n600), .A3(new_n671), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n664), .A2(new_n671), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n683), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n687), .A3(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n218), .B2(new_n693), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT28), .Z(new_n698));
  AND2_X1   g0498(.A1(new_n647), .A2(new_n645), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT26), .A3(new_n652), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT95), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n599), .A2(new_n552), .A3(new_n559), .A4(new_n647), .ZN(new_n703));
  AND4_X1   g0503(.A1(new_n602), .A2(new_n633), .A3(new_n636), .A4(new_n639), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n645), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n513), .A2(new_n518), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n652), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n654), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n701), .A3(new_n700), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n670), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n670), .B1(new_n651), .B2(new_n657), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(KEYINPUT96), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n711), .A2(new_n716), .A3(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n635), .A2(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n627), .A2(new_n520), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT87), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n627), .A2(new_n520), .A3(KEYINPUT87), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT93), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(G179), .A4(new_n626), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n489), .A2(new_n574), .A3(new_n495), .A4(new_n534), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(G179), .B1(new_n492), .B2(new_n493), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n535), .A2(new_n730), .A3(new_n571), .A4(new_n630), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT30), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT31), .A4(new_n670), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n671), .B1(new_n729), .B2(new_n732), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n737), .B2(new_n734), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT94), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n641), .A2(new_n671), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n733), .A2(new_n734), .A3(new_n670), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n735), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n718), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n698), .B1(new_n749), .B2(G1), .ZN(G364));
  NOR2_X1   g0550(.A1(new_n250), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n255), .B1(new_n751), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n693), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n678), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n676), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n214), .B1(G20), .B2(new_n319), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n692), .A2(new_n417), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G45), .B2(new_n217), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n248), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n291), .A2(new_n211), .ZN(new_n765));
  INV_X1    g0565(.A(G355), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n766), .B1(G116), .B2(new_n211), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n761), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n754), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n215), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n368), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n463), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n775), .A2(KEYINPUT32), .B1(new_n779), .B2(new_n205), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G87), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n215), .A2(new_n463), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT98), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n368), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n783), .B1(new_n789), .B2(new_n350), .C1(new_n202), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n770), .A2(new_n368), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n775), .A2(KEYINPUT32), .B1(G107), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n771), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n287), .B1(G77), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT97), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n784), .A2(new_n799), .A3(new_n776), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n784), .B2(new_n776), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n795), .B(new_n798), .C1(new_n802), .C2(new_n262), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G303), .B1(new_n790), .B2(G326), .ZN(new_n808));
  XOR2_X1   g0608(.A(KEYINPUT33), .B(G317), .Z(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n789), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n802), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G322), .ZN(new_n812));
  INV_X1    g0612(.A(new_n772), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n797), .B1(new_n813), .B2(G329), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n794), .A2(G283), .B1(new_n778), .B2(G294), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n812), .A2(new_n287), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n792), .A2(new_n803), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT100), .ZN(new_n818));
  INV_X1    g0618(.A(new_n760), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n817), .B2(KEYINPUT100), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n769), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n759), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n675), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n756), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  AOI21_X1  g0625(.A(new_n384), .B1(new_n813), .B2(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n350), .B2(new_n793), .C1(new_n262), .C2(new_n779), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n811), .A2(G143), .B1(G159), .B2(new_n797), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n789), .B2(new_n829), .C1(new_n830), .C2(new_n791), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT34), .Z(new_n832));
  AOI211_X1 g0632(.A(new_n827), .B(new_n832), .C1(G50), .C2(new_n807), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n834), .A2(new_n789), .B1(new_n791), .B2(new_n624), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n793), .A2(new_n221), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n287), .B1(new_n837), .B2(new_n772), .C1(new_n604), .C2(new_n796), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(G97), .C2(new_n778), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n802), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n835), .B(new_n841), .C1(G107), .C2(new_n807), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n760), .B1(new_n833), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n760), .A2(new_n757), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n843), .B(new_n754), .C1(G77), .C2(new_n845), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n462), .A2(new_n464), .A3(new_n670), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n670), .B1(new_n459), .B2(new_n461), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n469), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n466), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n846), .B1(new_n757), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n713), .B(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n747), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n754), .B1(new_n854), .B2(new_n747), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  OAI21_X1  g0659(.A(new_n544), .B1(new_n541), .B2(new_n545), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT35), .ZN(new_n861));
  OAI211_X1 g0661(.A(G116), .B(new_n216), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT36), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n218), .B(G77), .C1(new_n262), .C2(new_n350), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n202), .A2(G68), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n255), .B(G13), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n751), .A2(new_n255), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n442), .B1(new_n413), .B2(new_n428), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n413), .A2(new_n668), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n383), .A2(new_n388), .A3(new_n393), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n874), .B2(KEYINPUT101), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n395), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n427), .B1(new_n877), .B2(new_n376), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n442), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n442), .A2(KEYINPUT102), .A3(new_n878), .ZN(new_n882));
  INV_X1    g0682(.A(new_n668), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n877), .B2(new_n376), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n873), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n438), .B2(new_n446), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n870), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n884), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n447), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n884), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT102), .B1(new_n442), .B2(new_n878), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n434), .A2(new_n427), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n434), .A2(new_n883), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .A4(new_n442), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n655), .A2(new_n656), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n850), .B(new_n671), .C1(new_n901), .C2(new_n705), .ZN(new_n902));
  INV_X1    g0702(.A(new_n847), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n365), .A2(new_n670), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n904), .B(new_n371), .C1(new_n347), .C2(new_n365), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n365), .B(new_n670), .C1(new_n347), .C2(new_n371), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n902), .A2(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n437), .A2(new_n668), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT103), .A3(new_n897), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n872), .B1(new_n437), .B2(new_n445), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT103), .B1(new_n911), .B2(new_n897), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n870), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n899), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n888), .A2(new_n899), .A3(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n347), .A2(new_n365), .A3(new_n671), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n909), .B(new_n910), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n662), .A2(new_n321), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n718), .B2(new_n471), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n907), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n850), .B1(new_n927), .B2(new_n905), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT105), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n559), .A2(new_n552), .ZN(new_n930));
  AND4_X1   g0730(.A1(new_n633), .A2(new_n636), .A3(new_n638), .A4(new_n639), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n707), .A2(new_n683), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n743), .B1(new_n932), .B2(new_n670), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n735), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n737), .A2(KEYINPUT104), .A3(KEYINPUT31), .A4(new_n734), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n929), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n743), .A4(new_n740), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n928), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n917), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT40), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n888), .B2(new_n899), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n938), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n471), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(G330), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n869), .B1(new_n926), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n953), .A2(new_n954), .B1(new_n926), .B2(new_n952), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n868), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OR2_X1    g0757(.A1(new_n517), .A2(new_n671), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n699), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n645), .A2(new_n958), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n930), .B1(new_n558), .B2(new_n671), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n652), .A2(new_n670), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n683), .A3(new_n689), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n552), .B1(new_n968), .B2(new_n602), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n671), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n966), .A2(new_n967), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n964), .A2(new_n967), .A3(new_n965), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n970), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n686), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n749), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n690), .A2(new_n687), .A3(new_n970), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT45), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n970), .B1(new_n690), .B2(new_n687), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT44), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n686), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n686), .B1(new_n985), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n690), .B1(new_n685), .B2(new_n689), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n677), .B2(KEYINPUT109), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n677), .B(KEYINPUT109), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n991), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n983), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n693), .B(KEYINPUT41), .Z(new_n996));
  OAI21_X1  g0796(.A(new_n752), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n982), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n966), .A2(new_n759), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n779), .A2(new_n206), .B1(new_n793), .B2(new_n205), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n417), .B1(new_n813), .B2(G317), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n834), .B2(new_n796), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G303), .C2(new_n811), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G294), .A2(new_n788), .B1(new_n790), .B2(G311), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n807), .B2(G116), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n781), .A2(new_n604), .A3(KEYINPUT46), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1003), .B(new_n1004), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n291), .B1(new_n290), .B2(new_n793), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n790), .A2(G143), .B1(new_n1009), .B2(KEYINPUT110), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(KEYINPUT110), .B2(new_n1009), .C1(new_n773), .C2(new_n789), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n796), .A2(new_n202), .B1(new_n772), .B2(new_n830), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G68), .B2(new_n778), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n262), .B2(new_n781), .C1(new_n829), .C2(new_n802), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1008), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n760), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n762), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n761), .B1(new_n211), .B2(new_n455), .C1(new_n1019), .C2(new_n241), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n999), .A2(new_n754), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n998), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n994), .A2(new_n753), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n417), .B1(new_n813), .B2(G326), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n604), .B2(new_n793), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n811), .A2(G317), .B1(G303), .B2(new_n797), .ZN(new_n1026));
  INV_X1    g0826(.A(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n789), .B2(new_n837), .C1(new_n1027), .C2(new_n791), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n782), .A2(G294), .B1(new_n778), .B2(G283), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1025), .B1(new_n1035), .B2(KEYINPUT112), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT112), .B2(new_n1035), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G159), .A2(new_n790), .B1(new_n788), .B2(new_n266), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n290), .A2(new_n781), .B1(new_n793), .B2(new_n205), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n455), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n778), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n417), .B1(new_n772), .B2(new_n829), .C1(new_n350), .C2(new_n796), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n811), .B2(G50), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1038), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n819), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n762), .B1(new_n238), .B2(new_n299), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n695), .B2(new_n765), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n266), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n1048), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n1048), .B2(G50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n695), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1047), .A2(new_n1052), .B1(new_n206), .B2(new_n692), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n761), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n754), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n685), .B2(new_n822), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n994), .A2(new_n749), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n693), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n994), .A2(new_n749), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1023), .B(new_n1057), .C1(new_n1059), .C2(new_n1060), .ZN(G393));
  NAND2_X1  g0861(.A1(new_n990), .A2(new_n753), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n762), .A2(new_n245), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n761), .B1(new_n211), .B2(new_n205), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n754), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n790), .A2(G150), .B1(G159), .B2(new_n811), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n384), .B1(new_n813), .B2(G143), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1048), .B2(new_n796), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n779), .A2(new_n290), .B1(new_n793), .B2(new_n221), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G68), .C2(new_n782), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n202), .B2(new_n789), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n790), .A2(G317), .B1(G311), .B2(new_n811), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n206), .A2(new_n793), .B1(new_n781), .B2(new_n834), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n287), .B1(new_n840), .B2(new_n796), .C1(new_n1027), .C2(new_n772), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n608), .C2(new_n778), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n624), .B2(new_n789), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1067), .A2(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1065), .B1(new_n1079), .B2(new_n760), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n970), .B2(new_n822), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n990), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n693), .B1(new_n1082), .B2(new_n1058), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n990), .B1(new_n749), .B2(new_n994), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1062), .B(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(G390));
  OAI21_X1  g0885(.A(new_n754), .B1(new_n266), .B2(new_n845), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT116), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n779), .A2(new_n773), .B1(new_n793), .B2(new_n202), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n796), .A2(new_n1089), .B1(new_n772), .B2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1088), .A2(new_n1091), .A3(new_n287), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1092), .B1(new_n789), .B2(new_n830), .C1(new_n1093), .C2(new_n791), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n781), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT53), .B1(new_n781), .B2(new_n829), .ZN(new_n1096));
  INV_X1    g0896(.A(G132), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1096), .C1(new_n802), .C2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n807), .A2(G87), .B1(new_n788), .B2(G107), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n834), .B2(new_n791), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n811), .A2(G116), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G97), .A2(new_n797), .B1(new_n813), .B2(G294), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n794), .A2(G68), .B1(new_n778), .B2(G77), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n287), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1094), .A2(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1087), .B1(new_n1105), .B2(new_n760), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n919), .A2(new_n920), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n758), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n951), .B1(new_n940), .B2(new_n938), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n928), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT113), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n922), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n908), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n466), .A2(new_n849), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n847), .B1(new_n713), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n927), .A2(new_n905), .ZN(new_n1118));
  OAI211_X1 g0918(.A(KEYINPUT113), .B(new_n922), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n919), .B2(new_n920), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n706), .A2(new_n710), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n671), .A3(new_n1116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n903), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1126), .A2(new_n922), .A3(new_n917), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1112), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n748), .A2(new_n850), .A3(new_n1125), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n922), .A3(new_n917), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n1107), .C2(new_n1120), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1108), .B1(new_n1132), .B2(new_n752), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1135), .B(new_n1108), .C1(new_n1132), .C2(new_n752), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT115), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n471), .A2(new_n1109), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n925), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1109), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1118), .B1(new_n1141), .B2(new_n851), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1124), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1129), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1118), .B1(new_n747), .B2(new_n851), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1111), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1117), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT114), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT114), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1149), .B(new_n1117), .C1(new_n1111), .C2(new_n1145), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1144), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1137), .B1(new_n1140), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1132), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n693), .B1(new_n1152), .B2(new_n1132), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1134), .B(new_n1136), .C1(new_n1154), .C2(new_n1155), .ZN(G378));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n274), .A2(new_n883), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n318), .A2(new_n321), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n318), .B2(new_n321), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n946), .B2(G330), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT40), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n900), .A2(new_n941), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n917), .B2(new_n941), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n1166), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n923), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1166), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n942), .A2(KEYINPUT40), .B1(new_n941), .B2(new_n944), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n951), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n909), .A2(new_n910), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1178), .A3(new_n1171), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(KEYINPUT121), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1128), .A2(new_n1151), .A3(new_n1131), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1140), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT121), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1176), .A2(new_n1178), .A3(new_n1183), .A4(new_n1171), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT122), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1179), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1176), .A2(new_n1178), .A3(KEYINPUT122), .A4(new_n1171), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1173), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1186), .B1(new_n1181), .B2(new_n1140), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n694), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1180), .A2(new_n753), .A3(new_n1184), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n754), .B1(G50), .B2(new_n845), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n778), .A2(G150), .B1(new_n797), .B2(G137), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n781), .B2(new_n1089), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1090), .A2(new_n791), .B1(new_n789), .B2(new_n1097), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(G128), .C2(new_n811), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n773), .B2(new_n793), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT119), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n779), .A2(new_n350), .B1(new_n796), .B2(new_n455), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G107), .B2(new_n811), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n791), .B2(new_n614), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n384), .A2(new_n297), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G283), .B2(new_n813), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n262), .B2(new_n793), .C1(new_n290), .C2(new_n781), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT118), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1210), .B(new_n1214), .C1(G97), .C2(new_n788), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(KEYINPUT58), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1211), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1207), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1196), .B1(new_n1219), .B2(new_n760), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1166), .B2(new_n758), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT120), .Z(new_n1222));
  NAND2_X1  g1022(.A1(new_n1195), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1194), .A2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1140), .A2(new_n1151), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1149), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1146), .A2(KEYINPUT114), .A3(new_n1147), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1139), .A3(new_n1144), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n996), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1226), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1118), .A2(new_n757), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n754), .B1(G68), .B2(new_n845), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n807), .A2(G97), .B1(new_n788), .B2(new_n608), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n840), .B2(new_n791), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n811), .A2(G283), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G107), .A2(new_n797), .B1(new_n813), .B2(G303), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G77), .A2(new_n794), .B1(new_n778), .B2(new_n1040), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n287), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n790), .A2(G132), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n773), .B2(new_n806), .C1(new_n789), .C2(new_n1089), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n417), .B1(new_n796), .B2(new_n829), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G128), .B2(new_n813), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n794), .A2(G58), .B1(new_n778), .B2(G50), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n830), .C2(new_n802), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1237), .A2(new_n1241), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1235), .B1(new_n1248), .B2(new_n760), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1151), .A2(new_n753), .B1(new_n1234), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1233), .A2(new_n1250), .ZN(G381));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n858), .ZN(new_n1253));
  OR2_X1    g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1253), .A2(G387), .A3(new_n1254), .A4(G381), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1223), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1155), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1133), .B1(new_n1257), .B2(new_n1153), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .ZN(G407));
  NAND2_X1  g1059(.A1(new_n669), .A2(G213), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(G407), .A2(G213), .A3(new_n1262), .ZN(G409));
  XNOR2_X1  g1063(.A(G393), .B(new_n824), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n998), .A2(new_n1021), .A3(G390), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n998), .B2(new_n1021), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1252), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n998), .A2(new_n1021), .A3(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1264), .A3(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1268), .A2(new_n1271), .A3(KEYINPUT125), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT125), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1194), .A2(G378), .A3(new_n1224), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1191), .A2(new_n753), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1276), .B(new_n1222), .C1(new_n1185), .C2(new_n996), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1258), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1139), .A4(new_n1144), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n693), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1226), .A2(KEYINPUT60), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1231), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1250), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n858), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1231), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1280), .A2(new_n693), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(G384), .A3(new_n1250), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1279), .A2(new_n1260), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1261), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1261), .A2(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G384), .B1(new_n1288), .B2(new_n1250), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n858), .B(new_n1284), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1285), .A2(new_n1289), .A3(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1294), .B(new_n1295), .C1(new_n1296), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1296), .A2(new_n1305), .A3(new_n1291), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1293), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1256), .A2(G378), .B1(new_n1258), .B2(new_n1277), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1302), .B(new_n1301), .C1(new_n1308), .C2(new_n1261), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1294), .B1(new_n1309), .B2(new_n1295), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1274), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1309), .A2(KEYINPUT123), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1292), .A2(KEYINPUT63), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1296), .A2(new_n1314), .A3(new_n1291), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1268), .A2(new_n1271), .A3(new_n1295), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1309), .B2(KEYINPUT123), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1312), .A2(new_n1316), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1258), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1275), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1290), .A2(KEYINPUT126), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1258), .ZN(new_n1325));
  OAI221_X1 g1125(.A(new_n1275), .B1(new_n1256), .B2(new_n1325), .C1(KEYINPUT126), .C2(new_n1290), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1274), .A2(new_n1324), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1274), .A2(new_n1324), .A3(new_n1331), .A4(new_n1326), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1328), .A2(new_n1330), .A3(new_n1332), .ZN(G402));
endmodule


