//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n208), .B1(new_n209), .B2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT66), .B(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G58), .A2(G232), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n219), .B2(new_n222), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT70), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  INV_X1    g0049(.A(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT74), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G58), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n217), .A2(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n216), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(new_n271), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(G50), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  AND2_X1   g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n216), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(KEYINPUT72), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n291), .A2(new_n216), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n298), .A2(G1), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT71), .A2(G41), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT71), .A2(G41), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n304), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n271), .A2(new_n307), .B1(new_n293), .B2(new_n294), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n300), .A2(new_n305), .B1(G226), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n278), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n270), .A2(new_n275), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(KEYINPUT9), .B1(new_n256), .B2(KEYINPUT10), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n257), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n312), .A2(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(new_n257), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n316), .A4(new_n278), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n276), .C1(G169), .C2(new_n311), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n217), .ZN(new_n331));
  INV_X1    g0131(.A(new_n258), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n332), .A2(new_n202), .B1(new_n266), .B2(new_n286), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n269), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT11), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n330), .B2(new_n274), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n274), .A2(KEYINPUT12), .A3(G68), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(new_n272), .B2(G68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n300), .A2(new_n305), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n307), .A2(new_n271), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n293), .A2(new_n294), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n292), .A2(new_n295), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G226), .A2(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G232), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(G1698), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n283), .B1(G33), .B2(G97), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n344), .B1(new_n224), .B2(new_n347), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n352), .A2(new_n348), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n308), .A2(G238), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n344), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n358), .A3(KEYINPUT75), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(new_n360), .A3(KEYINPUT13), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(G169), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g0163(.A(new_n358), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n322), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n362), .A2(KEYINPUT14), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n343), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n342), .B1(new_n370), .B2(new_n354), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n359), .A2(G200), .A3(new_n361), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(KEYINPUT77), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G20), .A2(G77), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n378), .B1(new_n260), .B2(new_n332), .C1(new_n266), .C2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n380), .A2(new_n269), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n272), .A2(G77), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G77), .B2(new_n274), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G244), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n344), .B1(new_n385), .B2(new_n347), .ZN(new_n386));
  AND2_X1   g0186(.A1(KEYINPUT3), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(KEYINPUT3), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G107), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n283), .A2(new_n284), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n391), .B2(new_n350), .C1(new_n224), .C2(new_n287), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n392), .B2(new_n296), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G169), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n384), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n322), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n394), .A2(G200), .ZN(new_n400));
  INV_X1    g0200(.A(new_n384), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(G190), .B2(new_n393), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n326), .A2(new_n368), .A3(new_n377), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT80), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n265), .A2(new_n272), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n274), .B2(new_n265), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n281), .A2(new_n217), .A3(new_n282), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n282), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n413), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n330), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n220), .B1(new_n223), .B2(new_n263), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n269), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n258), .A2(G159), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n201), .B1(new_n330), .B2(G58), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n217), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n250), .B1(new_n411), .B2(new_n413), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n423), .B1(new_n428), .B2(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n408), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n300), .A2(new_n305), .B1(G232), .B2(new_n308), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n288), .A2(new_n284), .ZN(new_n432));
  INV_X1    g0232(.A(G226), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G1698), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n432), .B(new_n434), .C1(new_n387), .C2(new_n388), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n296), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n431), .A2(G179), .A3(new_n438), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT18), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n408), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT7), .B1(new_n389), .B2(new_n217), .ZN(new_n446));
  OAI21_X1  g0246(.A(G68), .B1(new_n446), .B2(new_n415), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n419), .A2(new_n447), .A3(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n269), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT16), .B1(new_n417), .B2(new_n419), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n442), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n348), .B1(new_n436), .B2(new_n435), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT71), .B(G41), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G45), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n346), .A2(new_n271), .A3(G274), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n457), .A2(new_n458), .B1(new_n347), .B2(new_n350), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n455), .A2(new_n459), .A3(new_n369), .ZN(new_n460));
  INV_X1    g0260(.A(G200), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n431), .B2(new_n438), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n454), .B1(new_n451), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n422), .A2(new_n429), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n460), .A2(new_n462), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(KEYINPUT17), .A3(new_n445), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n444), .A2(new_n453), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  XOR2_X1   g0268(.A(new_n468), .B(KEYINPUT79), .Z(new_n469));
  NAND3_X1  g0269(.A1(new_n405), .A2(new_n406), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT80), .B1(new_n471), .B2(new_n404), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n414), .A2(G107), .A3(new_n416), .ZN(new_n474));
  INV_X1    g0274(.A(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  XOR2_X1   g0276(.A(G97), .B(G107), .Z(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n423), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n271), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n423), .A2(new_n274), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G97), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G97), .B2(new_n274), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n480), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT5), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n301), .B2(new_n302), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n304), .A2(G1), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n346), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  INV_X1    g0300(.A(new_n498), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n298), .A2(new_n299), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n496), .A4(new_n495), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n500), .B1(new_n499), .B2(new_n503), .ZN(new_n506));
  OAI211_X1 g0306(.A(G250), .B(G1698), .C1(new_n387), .C2(new_n388), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n283), .A2(G244), .A3(new_n284), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(KEYINPUT4), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n348), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR4_X1   g0315(.A1(new_n505), .A2(new_n506), .A3(new_n322), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n499), .A2(new_n503), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(KEYINPUT82), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n395), .B1(new_n518), .B2(new_n504), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n490), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(G190), .A3(new_n504), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n505), .A2(new_n506), .A3(new_n515), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n486), .C1(new_n522), .C2(new_n461), .ZN(new_n523));
  NAND3_X1  g0323(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n217), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n206), .B2(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n217), .B(G68), .C1(new_n387), .C2(new_n388), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n266), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT84), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n526), .A2(new_n533), .A3(new_n527), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n269), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n379), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n483), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n274), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n379), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G238), .B(new_n284), .C1(new_n387), .C2(new_n388), .ZN(new_n541));
  OAI211_X1 g0341(.A(G244), .B(G1698), .C1(new_n387), .C2(new_n388), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n296), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n494), .A2(new_n299), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n546), .B(new_n346), .C1(G250), .C2(new_n494), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n322), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n547), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n395), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(G190), .A3(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(G200), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n535), .A2(new_n539), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n483), .A2(G87), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n549), .A2(new_n551), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n520), .A2(new_n523), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n217), .B(G87), .C1(new_n387), .C2(new_n388), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n283), .A2(new_n563), .A3(new_n217), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n543), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n217), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n475), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n566), .B1(new_n565), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n269), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G264), .B(new_n346), .C1(new_n497), .C2(new_n498), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n391), .A2(new_n576), .B1(new_n280), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n296), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n575), .A2(new_n581), .A3(new_n503), .A4(G190), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n538), .A2(new_n475), .ZN(new_n583));
  NOR2_X1   g0383(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n585), .A2(new_n587), .B1(new_n483), .B2(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n574), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(new_n581), .A3(new_n503), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n574), .A2(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n395), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(G179), .C2(new_n590), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G116), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n268), .A2(new_n216), .B1(G20), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n508), .B(new_n217), .C1(G33), .C2(new_n529), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(KEYINPUT85), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n538), .A2(new_n597), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n482), .C2(new_n597), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n600), .A2(KEYINPUT85), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n600), .A2(KEYINPUT85), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n598), .C2(new_n599), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G270), .B(new_n346), .C1(new_n497), .C2(new_n498), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n283), .A2(G257), .A3(new_n284), .ZN(new_n610));
  INV_X1    g0410(.A(G303), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n283), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n296), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n503), .A3(new_n613), .A4(G190), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n503), .A3(new_n613), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n607), .B(new_n614), .C1(new_n616), .C2(new_n461), .ZN(new_n617));
  INV_X1    g0417(.A(new_n607), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n618), .A3(G169), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n503), .A2(new_n613), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n618), .A3(G179), .A4(new_n608), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n615), .A2(new_n618), .A3(KEYINPUT21), .A4(G169), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n617), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n623), .A2(new_n624), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT86), .A3(new_n621), .A4(new_n617), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n596), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n473), .A2(new_n560), .A3(new_n630), .ZN(G372));
  NOR2_X1   g0431(.A1(new_n589), .A2(new_n591), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n540), .A2(new_n548), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n545), .A2(KEYINPUT88), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n544), .A2(new_n296), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n547), .B(KEYINPUT89), .Z(new_n638));
  AOI21_X1  g0438(.A(G169), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n461), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n535), .A2(new_n552), .A3(new_n539), .A4(new_n556), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n633), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n520), .A2(new_n643), .A3(new_n523), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT90), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n520), .A2(new_n643), .A3(new_n523), .A4(KEYINPUT90), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n628), .A2(new_n595), .A3(new_n621), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n559), .B(new_n490), .C1(new_n516), .C2(new_n519), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n517), .A2(KEYINPUT82), .ZN(new_n652));
  INV_X1    g0452(.A(new_n515), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n504), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G169), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n322), .B2(new_n654), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n642), .ZN(new_n658));
  INV_X1    g0458(.A(new_n486), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n639), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n549), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n651), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n649), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n473), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n324), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n451), .A2(new_n452), .A3(new_n442), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n452), .B1(new_n451), .B2(new_n442), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n367), .B1(new_n377), .B2(new_n399), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n464), .A2(new_n467), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n318), .A2(new_n321), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n665), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n271), .A2(new_n217), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n607), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n627), .B2(new_n629), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n628), .A2(new_n621), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n683), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n593), .A2(new_n681), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n592), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(new_n595), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n595), .A2(new_n681), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n685), .A2(new_n682), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n213), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n456), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n703), .A2(new_n271), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n221), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n703), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n637), .A2(new_n638), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n322), .A3(new_n615), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n654), .A2(new_n590), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(KEYINPUT91), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n654), .A2(new_n715), .A3(new_n590), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n575), .A2(new_n581), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n550), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n616), .A2(new_n717), .A3(G179), .A4(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT92), .B(KEYINPUT30), .C1(new_n721), .C2(new_n654), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n615), .A2(new_n322), .ZN(new_n723));
  NAND2_X1  g0523(.A1(KEYINPUT92), .A2(KEYINPUT30), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n717), .A2(new_n720), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n522), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n714), .A2(new_n716), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n682), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n710), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n590), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT91), .B1(new_n522), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n712), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n716), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n722), .A2(new_n726), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT93), .A3(new_n729), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n682), .B1(new_n735), .B2(new_n736), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n520), .A2(new_n523), .A3(new_n559), .A4(new_n682), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n742), .A2(new_n728), .B1(new_n744), .B2(new_n630), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n689), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n681), .B1(new_n649), .B2(new_n663), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n656), .A2(new_n659), .A3(new_n658), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT26), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n520), .A2(new_n648), .A3(new_n643), .A4(new_n523), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n749), .A2(new_n751), .A3(new_n662), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .A3(new_n682), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n746), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n709), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n211), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n271), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n703), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n216), .B1(G20), .B2(new_n395), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n217), .A2(new_n322), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n389), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n217), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n765), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n768), .B1(G329), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n764), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n369), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n322), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(G294), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n764), .A2(new_n776), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT95), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n780), .B1(G322), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n773), .A2(new_n369), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n769), .A2(new_n369), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n789), .A2(G326), .B1(new_n791), .B2(G283), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n788), .B(new_n792), .C1(new_n611), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n789), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT96), .B(G159), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n771), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n795), .A2(new_n202), .B1(new_n798), .B2(KEYINPUT32), .ZN(new_n799));
  INV_X1    g0599(.A(new_n774), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n800), .A2(new_n250), .B1(new_n790), .B2(new_n475), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n787), .A2(G58), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n283), .B1(new_n766), .B2(new_n286), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n798), .B2(KEYINPUT32), .ZN(new_n805));
  INV_X1    g0605(.A(new_n793), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G87), .B1(new_n778), .B2(G97), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n763), .B1(new_n794), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n762), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n213), .A2(G355), .A3(new_n283), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n702), .A2(new_n283), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n222), .B2(G45), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n254), .A2(new_n304), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n814), .B1(G116), .B2(new_n213), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n761), .B(new_n809), .C1(new_n813), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n688), .ZN(new_n820));
  INV_X1    g0620(.A(new_n812), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n688), .A2(new_n689), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT94), .ZN(new_n824));
  INV_X1    g0624(.A(new_n690), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n761), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(G396));
  INV_X1    g0627(.A(new_n747), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n402), .A2(new_n400), .B1(new_n401), .B2(new_n681), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n399), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n398), .A2(new_n681), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n833), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n664), .A2(new_n682), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n746), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n760), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n835), .A2(new_n746), .A3(new_n837), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n762), .A2(new_n810), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n761), .B1(new_n286), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(KEYINPUT97), .B(G283), .Z(new_n844));
  OAI22_X1  g0644(.A1(new_n800), .A2(new_n844), .B1(new_n793), .B2(new_n475), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n389), .B1(new_n766), .B2(new_n597), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G311), .B2(new_n771), .ZN(new_n847));
  INV_X1    g0647(.A(G87), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n790), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G97), .B2(new_n778), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n847), .B(new_n850), .C1(new_n786), .C2(new_n577), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n845), .B(new_n851), .C1(G303), .C2(new_n789), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n283), .B1(new_n770), .B2(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n202), .A2(new_n793), .B1(new_n790), .B2(new_n250), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(G58), .C2(new_n778), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT98), .Z(new_n857));
  INV_X1    g0657(.A(new_n766), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n789), .A2(G137), .B1(new_n797), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n859), .B1(new_n860), .B2(new_n800), .C1(new_n786), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n852), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n843), .B1(new_n763), .B2(new_n864), .C1(new_n836), .C2(new_n811), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n841), .A2(new_n865), .ZN(G384));
  XOR2_X1   g0666(.A(new_n478), .B(KEYINPUT100), .Z(new_n867));
  INV_X1    g0667(.A(KEYINPUT35), .ZN(new_n868));
  OAI211_X1 g0668(.A(G116), .B(new_n218), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n707), .B(G77), .C1(new_n263), .C2(new_n223), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n271), .B(G13), .C1(new_n872), .C2(new_n249), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n451), .A2(new_n442), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n466), .B(new_n445), .C1(new_n450), .C2(new_n449), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  INV_X1    g0679(.A(new_n679), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n451), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(KEYINPUT103), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n876), .A2(new_n881), .A3(new_n877), .A4(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n448), .A3(new_n269), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n445), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n445), .A3(KEYINPUT102), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n880), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n442), .A3(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n877), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n882), .A2(new_n885), .B1(KEYINPUT37), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n671), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n896), .B2(new_n669), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n875), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n897), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n883), .B(KEYINPUT103), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(KEYINPUT38), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT39), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n367), .A2(new_n682), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n882), .A2(new_n885), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT105), .A3(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n881), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n468), .A2(KEYINPUT104), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT104), .B1(new_n468), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n878), .A2(new_n881), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n907), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n904), .B(new_n906), .C1(new_n921), .C2(KEYINPUT39), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n679), .B1(new_n667), .B2(new_n668), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n898), .A2(new_n902), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n343), .A2(new_n682), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n375), .A2(new_n376), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n367), .ZN(new_n927));
  INV_X1    g0727(.A(new_n925), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n368), .A2(new_n377), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n837), .B2(new_n832), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT101), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n831), .B1(new_n747), .B2(new_n836), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n935), .A2(KEYINPUT101), .A3(new_n931), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n922), .B(new_n923), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n473), .A2(new_n748), .A3(new_n754), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n674), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n833), .B1(new_n927), .B2(new_n929), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n744), .A2(new_n630), .B1(new_n737), .B2(new_n729), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT106), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT106), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n944), .B(new_n728), .C1(new_n727), .C2(new_n682), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT40), .B1(new_n921), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n941), .A2(new_n946), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT40), .B1(new_n898), .B2(new_n902), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n473), .A2(new_n946), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n689), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n940), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n271), .B2(new_n757), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n940), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n874), .B1(new_n957), .B2(new_n958), .ZN(G367));
  INV_X1    g0759(.A(new_n695), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n520), .B(new_n523), .C1(new_n486), .C2(new_n682), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n656), .A2(new_n659), .A3(new_n681), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n960), .A2(new_n964), .A3(new_n698), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n520), .B1(new_n964), .B2(new_n595), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n682), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n681), .B1(new_n555), .B2(new_n557), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n658), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n662), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n966), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n972), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n696), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n966), .A2(new_n975), .A3(new_n974), .A4(new_n968), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n963), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n696), .B2(new_n964), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n703), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n964), .A2(new_n699), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT44), .Z(new_n987));
  AND3_X1   g0787(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT45), .B1(new_n700), .B2(new_n963), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(KEYINPUT108), .A3(new_n978), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n695), .B(new_n698), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n825), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n755), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n978), .A2(KEYINPUT108), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n985), .B1(new_n998), .B2(new_n755), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n980), .B(new_n982), .C1(new_n999), .C2(new_n759), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n815), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n244), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n813), .B1(new_n213), .B2(new_n379), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n760), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n786), .A2(new_n860), .ZN(new_n1005));
  INV_X1    g0805(.A(G137), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n283), .B1(new_n770), .B2(new_n1006), .C1(new_n202), .C2(new_n766), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n800), .A2(new_n796), .B1(new_n790), .B2(new_n286), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n778), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n250), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G143), .B2(new_n789), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n263), .C2(new_n793), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n800), .A2(new_n577), .B1(new_n790), .B2(new_n529), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n786), .A2(new_n611), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n795), .A2(new_n767), .B1(new_n1010), .B2(new_n475), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n389), .B1(new_n770), .B2(new_n1017), .C1(new_n844), .C2(new_n766), .ZN(new_n1018));
  OR4_X1    g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT109), .B1(new_n806), .B2(G116), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT46), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n1013), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1004), .B1(new_n1023), .B2(new_n762), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n821), .B2(new_n972), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1000), .A2(new_n1025), .ZN(G387));
  NAND3_X1  g0826(.A1(new_n705), .A2(new_n213), .A3(new_n283), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(G107), .B2(new_n213), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n240), .A2(new_n304), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT110), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n304), .B1(new_n250), .B2(new_n286), .C1(new_n705), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n705), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n260), .A2(G50), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1001), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1028), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n813), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n760), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n774), .A2(G311), .B1(new_n858), .B2(G303), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n795), .C1(new_n786), .C2(new_n1017), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1010), .A2(new_n844), .B1(new_n793), .B2(new_n577), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n790), .A2(new_n597), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n283), .B(new_n1050), .C1(G326), .C2(new_n771), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n787), .A2(G50), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n806), .A2(G77), .B1(new_n791), .B2(G97), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n283), .B1(new_n770), .B2(new_n860), .C1(new_n250), .C2(new_n766), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n265), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n774), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n789), .A2(G159), .B1(new_n778), .B2(new_n536), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n763), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1038), .B(new_n1060), .C1(new_n960), .C2(new_n812), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n993), .B2(new_n759), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n994), .A2(new_n703), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n755), .A2(new_n993), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(G393));
  NAND2_X1  g0865(.A1(new_n990), .A2(new_n978), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n987), .B(new_n696), .C1(new_n988), .C2(new_n989), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n759), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1001), .A2(new_n248), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n813), .B1(new_n529), .B2(new_n213), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n760), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n786), .A2(new_n767), .B1(new_n1017), .B2(new_n795), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT52), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n800), .A2(new_n611), .B1(new_n790), .B2(new_n475), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1010), .A2(new_n597), .B1(new_n844), .B2(new_n793), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n389), .B1(new_n770), .B2(new_n1040), .C1(new_n577), .C2(new_n766), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n787), .A2(G159), .B1(G150), .B2(new_n789), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n800), .A2(new_n202), .B1(new_n223), .B2(new_n793), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1010), .A2(new_n286), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n283), .B1(new_n770), .B2(new_n861), .C1(new_n260), .C2(new_n766), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n849), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1073), .A2(new_n1077), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1071), .B1(new_n1087), .B2(new_n762), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n963), .B2(new_n821), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1068), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT112), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT112), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1068), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n998), .A2(new_n703), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n994), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1098), .ZN(G390));
  NAND3_X1  g0899(.A1(new_n746), .A2(new_n836), .A3(new_n930), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n946), .A2(G330), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n931), .B1(new_n1101), .B2(new_n834), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n753), .A2(new_n682), .A3(new_n830), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n832), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT113), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n627), .A2(new_n629), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n596), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1110), .A2(new_n743), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n836), .C1(new_n739), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n931), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n941), .A2(new_n946), .A3(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n837), .A2(new_n832), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(KEYINPUT113), .B(new_n935), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1106), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n946), .A2(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n473), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n938), .A2(new_n674), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1104), .A2(new_n930), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n895), .A2(new_n911), .A3(new_n897), .A4(new_n875), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT105), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n468), .A2(new_n913), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT104), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n468), .A2(KEYINPUT104), .A3(new_n913), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n882), .A2(new_n885), .B1(new_n917), .B2(KEYINPUT37), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n875), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1126), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1125), .A2(new_n905), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n906), .B1(new_n1116), .B2(new_n930), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT39), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n924), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1100), .B(new_n1136), .C1(new_n1137), .C2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n904), .B1(new_n921), .B2(KEYINPUT39), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n905), .B1(new_n935), .B2(new_n931), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n905), .B(new_n910), .C1(new_n912), .C2(new_n920), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1142), .A2(new_n1143), .B1(new_n1145), .B2(new_n1125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1141), .B1(new_n1146), .B2(new_n1114), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1124), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n703), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1124), .B2(new_n1147), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1142), .A2(new_n810), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1082), .B1(new_n787), .B2(G116), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT116), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n389), .B1(new_n770), .B2(new_n577), .C1(new_n529), .C2(new_n766), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n250), .A2(new_n790), .B1(new_n793), .B2(new_n848), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n789), .A2(G283), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n800), .B2(new_n475), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n283), .B1(new_n790), .B2(new_n202), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT115), .Z(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n766), .A2(new_n1162), .B1(new_n770), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1165), .A2(new_n795), .B1(new_n800), .B2(new_n1006), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G159), .C2(new_n778), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT53), .B1(new_n793), .B2(new_n860), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n793), .A2(KEYINPUT53), .A3(new_n860), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n787), .B2(G132), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1161), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n762), .B1(new_n1159), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n761), .B1(new_n265), .B2(new_n842), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT114), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1152), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT117), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1152), .A2(KEYINPUT117), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1141), .B(new_n759), .C1(new_n1146), .C2(new_n1114), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(KEYINPUT118), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT118), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1151), .B1(new_n1182), .B2(new_n1183), .ZN(G378));
  NOR2_X1   g0984(.A1(new_n315), .A2(new_n679), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n325), .B(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n952), .B2(G330), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n689), .B(new_n1188), .C1(new_n948), .C2(new_n951), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n937), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n910), .A3(new_n946), .A4(new_n941), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1194), .A2(KEYINPUT40), .B1(new_n949), .B2(new_n950), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1195), .B2(new_n689), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1116), .A2(new_n930), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n903), .B1(new_n1197), .B2(KEYINPUT101), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n936), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n922), .A2(new_n923), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT40), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n949), .B2(new_n1135), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n947), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G330), .B(new_n1189), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1196), .A2(new_n1200), .A3(new_n1202), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1192), .A2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1100), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1120), .A2(new_n941), .B1(new_n1112), .B2(new_n931), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT113), .B1(new_n1210), .B2(new_n935), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1115), .A2(new_n1107), .A3(new_n1116), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1209), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1123), .B1(new_n1147), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1208), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT57), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT119), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1192), .A2(new_n1207), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n937), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1220), .A2(KEYINPUT119), .A3(new_n1196), .A4(new_n1206), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1214), .A4(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1217), .A2(new_n703), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G33), .A2(G41), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G50), .B(new_n1224), .C1(new_n303), .C2(new_n389), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n456), .B(new_n283), .C1(new_n771), .C2(G283), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n379), .B2(new_n766), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1011), .B(new_n1227), .C1(G77), .C2(new_n806), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n529), .A2(new_n800), .B1(new_n795), .B2(new_n597), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G58), .B2(new_n791), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n475), .C2(new_n786), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT58), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n800), .A2(new_n853), .B1(new_n766), .B2(new_n1006), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n787), .B2(G128), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n789), .A2(G125), .B1(new_n778), .B2(G150), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n793), .C2(new_n1162), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1240));
  INV_X1    g1040(.A(G124), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1224), .B1(new_n770), .B2(new_n1241), .C1(new_n796), .C2(new_n790), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n762), .B1(new_n1234), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n761), .B1(new_n202), .B2(new_n842), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n1189), .C2(new_n811), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1208), .B2(new_n759), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1223), .A2(new_n1248), .ZN(G375));
  OAI211_X1 g1049(.A(new_n1122), .B(new_n1106), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1124), .A2(new_n984), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n931), .A2(new_n810), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT120), .ZN(new_n1253));
  INV_X1    g1053(.A(G159), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n793), .A2(new_n1254), .B1(new_n770), .B2(new_n1165), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n853), .A2(new_n795), .B1(new_n800), .B2(new_n1162), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(G137), .C2(new_n787), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n283), .B1(new_n790), .B2(new_n263), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT122), .Z(new_n1259));
  AOI22_X1  g1059(.A1(G50), .A2(new_n778), .B1(new_n858), .B2(G150), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT121), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n800), .A2(new_n597), .B1(new_n793), .B2(new_n529), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G294), .B2(new_n789), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n787), .A2(G283), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n389), .B1(new_n770), .B2(new_n611), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G107), .B2(new_n858), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G77), .A2(new_n791), .B1(new_n778), .B2(new_n536), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1264), .A2(new_n1265), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n763), .B1(new_n1262), .B2(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n761), .B(new_n1270), .C1(new_n250), .C2(new_n842), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1119), .A2(new_n759), .B1(new_n1253), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1251), .A2(new_n1272), .ZN(G381));
  NOR4_X1   g1073(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1000), .A3(new_n1025), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G378), .A2(new_n1275), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1076(.A(new_n1183), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1277), .A2(new_n1181), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G213), .A3(new_n680), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(G375), .C2(new_n1279), .ZN(G409));
  NAND3_X1  g1080(.A1(new_n1223), .A2(G378), .A3(new_n1248), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1219), .A2(new_n759), .A3(new_n1221), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1246), .C1(new_n985), .C2(new_n1215), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1278), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n680), .A2(G213), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1149), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1213), .A2(KEYINPUT60), .A3(new_n1122), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1250), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT123), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT123), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .A4(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1295));
  AND4_X1   g1095(.A1(new_n1272), .A2(new_n1292), .A3(new_n1294), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1272), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1291), .B2(KEYINPUT123), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1301), .B2(new_n1294), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1285), .A2(new_n1286), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1292), .A2(new_n1272), .A3(new_n1294), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1298), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1301), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n680), .A2(G213), .A3(G2897), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1310), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1306), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1281), .A2(new_n1284), .B1(G213), .B2(new_n680), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1303), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1305), .A2(new_n1314), .A3(new_n1315), .A4(new_n1318), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1093), .A2(new_n1091), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G390), .A2(new_n1000), .A3(new_n1025), .ZN(new_n1322));
  XOR2_X1   g1122(.A(G393), .B(G396), .Z(new_n1323));
  AND3_X1   g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1313), .A2(new_n1311), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1315), .B(new_n1326), .C1(new_n1329), .C2(new_n1316), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1304), .A2(KEYINPUT125), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1304), .A2(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT63), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1331), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1328), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1278), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1303), .ZN(new_n1341));
  OAI211_X1 g1141(.A(G375), .B(new_n1278), .C1(new_n1296), .C2(new_n1302), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1339), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(new_n1339), .A3(new_n1342), .ZN(new_n1346));
  OR3_X1    g1146(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT127), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .A4(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1346), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1327), .B(KEYINPUT127), .C1(new_n1349), .C2(new_n1343), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(G402));
endmodule


