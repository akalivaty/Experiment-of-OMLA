//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n210), .B1(new_n217), .B2(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n219), .A3(new_n216), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(KEYINPUT15), .A3(new_n210), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(KEYINPUT17), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n225), .B1(new_n221), .B2(new_n222), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n209), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n223), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n208), .B(new_n223), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n228), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n228), .A4(new_n229), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G169gat), .B(G197gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT12), .Z(new_n242));
  NAND4_X1  g041(.A1(new_n232), .A2(new_n235), .A3(new_n236), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT86), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n236), .A2(new_n235), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n232), .A4(new_n242), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n232), .ZN(new_n249));
  INV_X1    g048(.A(new_n242), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G8gat), .B(G36gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT75), .ZN(new_n255));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260));
  INV_X1    g059(.A(G211gat), .ZN(new_n261));
  INV_X1    g060(.A(G218gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n270));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n271), .C1(new_n272), .C2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n276), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT68), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n294), .B(KEYINPUT67), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n291), .B1(new_n287), .B2(new_n289), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n299), .C1(new_n285), .C2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n269), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n275), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT23), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n297), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n285), .B1(new_n292), .B2(KEYINPUT24), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT65), .B(G176gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g115(.A(new_n268), .B(new_n284), .C1(new_n307), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n284), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n307), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n307), .B2(new_n316), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n323));
  INV_X1    g122(.A(new_n268), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n267), .B(new_n317), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n324), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n284), .B1(new_n307), .B2(new_n316), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n266), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n258), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n267), .ZN(new_n334));
  INV_X1    g133(.A(new_n317), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n307), .A2(new_n316), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n307), .A2(new_n319), .A3(new_n316), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n284), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n325), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n335), .B(new_n266), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n341), .A3(new_n257), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(KEYINPUT30), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n334), .A2(new_n344), .A3(new_n341), .A4(new_n257), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT0), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT1), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G113gat), .A2(G120gat), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G127gat), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G134gat), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n355), .ZN(new_n366));
  AND4_X1   g165(.A1(new_n365), .A2(new_n366), .A3(new_n359), .A4(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G113gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n364), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n354), .B1(new_n368), .B2(new_n370), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT72), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n363), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT77), .B1(new_n383), .B2(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G148gat), .ZN(new_n387));
  INV_X1    g186(.A(G148gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G141gat), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n387), .A2(new_n389), .B1(KEYINPUT2), .B2(new_n381), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n377), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n364), .A3(new_n372), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT72), .B1(new_n374), .B2(new_n375), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n362), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(KEYINPUT2), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n388), .A2(G141gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n386), .A2(G148gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n384), .B2(new_n382), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n395), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n353), .B1(new_n398), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n377), .B2(new_n397), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n396), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n377), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n408), .A3(KEYINPUT4), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(new_n417), .A3(new_n352), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n353), .C1(new_n398), .C2(new_n409), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n419), .A2(KEYINPUT5), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n347), .B(new_n351), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(new_n351), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT6), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n351), .A3(new_n423), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT79), .B1(new_n346), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n266), .A2(new_n323), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n415), .B1(new_n432), .B2(KEYINPUT81), .ZN(new_n433));
  INV_X1    g232(.A(new_n323), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n267), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n397), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n266), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n431), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n415), .B1(new_n266), .B2(KEYINPUT29), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n397), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n441), .A2(new_n438), .A3(new_n431), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n439), .A2(G22gat), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT31), .B(G50gat), .Z(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT80), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(G22gat), .B1(new_n439), .B2(new_n442), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n443), .A2(new_n453), .A3(new_n450), .A4(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n427), .A2(new_n428), .ZN(new_n456));
  INV_X1    g255(.A(new_n424), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n343), .A2(new_n345), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n430), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n353), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n398), .A2(new_n409), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n464), .B(KEYINPUT39), .C1(new_n353), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n467), .A3(new_n353), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n468), .A2(new_n469), .A3(new_n351), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n468), .B2(new_n351), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n425), .A2(new_n426), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT40), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(new_n459), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n258), .A2(KEYINPUT37), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n332), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n334), .A2(new_n341), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n258), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n335), .B(new_n267), .C1(new_n339), .C2(new_n340), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n267), .B1(new_n327), .B2(new_n330), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n479), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n342), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n475), .A2(new_n492), .A3(new_n347), .A4(new_n428), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n457), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n427), .B2(new_n428), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n478), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n462), .B1(new_n497), .B2(new_n455), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n322), .A2(new_n401), .ZN(new_n499));
  INV_X1    g298(.A(G227gat), .ZN(new_n500));
  INV_X1    g299(.A(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n377), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT32), .ZN(new_n505));
  XOR2_X1   g304(.A(G15gat), .B(G43gat), .Z(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G99gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(new_n503), .ZN(new_n513));
  INV_X1    g312(.A(new_n502), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT34), .B(new_n502), .C1(new_n499), .C2(new_n503), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n505), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n508), .ZN(new_n522));
  INV_X1    g321(.A(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n513), .A2(new_n514), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT34), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n505), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n517), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n520), .B(new_n528), .C1(new_n529), .C2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n526), .A2(new_n527), .A3(new_n517), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n527), .B1(new_n526), .B2(new_n517), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n534), .A2(new_n535), .B1(new_n530), .B2(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n498), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n430), .A2(new_n461), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n444), .A2(new_n448), .B1(new_n443), .B2(new_n450), .ZN(new_n540));
  INV_X1    g339(.A(new_n454), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n528), .A3(new_n520), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT35), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n496), .A2(KEYINPUT35), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n534), .A2(new_n535), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n542), .A3(new_n546), .A4(new_n459), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n253), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(G57gat), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g354(.A1(new_n551), .A2(new_n552), .B1(new_n555), .B2(KEYINPUT9), .ZN(new_n556));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n209), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n209), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT88), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G155gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n575), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G127gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n360), .ZN(new_n581));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n579), .B2(new_n581), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n572), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(new_n584), .A3(new_n571), .A4(new_n569), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591));
  AND2_X1   g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT91), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(G85gat), .A3(G92gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(KEYINPUT7), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  OAI211_X1 g399(.A(KEYINPUT91), .B(new_n600), .C1(new_n594), .C2(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n594), .B2(new_n595), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n607), .A2(new_n599), .A3(new_n601), .A4(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n593), .B1(new_n610), .B2(new_n223), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT92), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n221), .B2(new_n222), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n593), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n609), .B1(new_n224), .B2(new_n226), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n591), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT93), .ZN(new_n624));
  INV_X1    g423(.A(new_n591), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT90), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n622), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n622), .B2(new_n626), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n590), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n590), .B(KEYINPUT94), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n608), .B(new_n606), .C1(new_n573), .C2(KEYINPUT95), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n608), .A2(KEYINPUT95), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n609), .A2(new_n559), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n559), .ZN(new_n642));
  INV_X1    g441(.A(G230gat), .ZN(new_n643));
  OAI22_X1  g442(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n501), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n501), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n638), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n646), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n549), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n458), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n459), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G8gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  MUX2_X1   g462(.A(new_n661), .B(new_n663), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g463(.A1(new_n532), .A2(new_n529), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n534), .A2(new_n535), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n532), .B1(new_n520), .B2(new_n528), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT96), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n533), .A2(new_n536), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n675), .B2(new_n656), .ZN(new_n676));
  INV_X1    g475(.A(new_n546), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n656), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT98), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n549), .A2(new_n455), .A3(new_n655), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  NAND3_X1  g484(.A1(new_n498), .A2(new_n668), .A3(new_n670), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n548), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n631), .A2(new_n632), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n538), .A2(new_n548), .ZN(new_n691));
  INV_X1    g490(.A(new_n688), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n690), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n253), .A2(new_n654), .A3(new_n590), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n458), .ZN(new_n701));
  INV_X1    g500(.A(new_n654), .ZN(new_n702));
  INV_X1    g501(.A(new_n590), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n549), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G29gat), .A3(new_n458), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n701), .A2(new_n708), .ZN(G1328gat));
  OAI21_X1  g508(.A(G36gat), .B1(new_n700), .B2(new_n459), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n706), .A2(G36gat), .A3(new_n459), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1329gat));
  OAI21_X1  g512(.A(G43gat), .B1(new_n696), .B2(new_n671), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n677), .A2(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT103), .B1(new_n706), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(KEYINPUT47), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n697), .A2(new_n674), .A3(new_n699), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(G43gat), .B1(new_n718), .B2(new_n717), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n722), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g522(.A1(new_n542), .A2(G50gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT105), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n726), .A2(KEYINPUT48), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT106), .B1(new_n696), .B2(new_n542), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n542), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n725), .B(KEYINPUT104), .Z(new_n733));
  NAND3_X1  g532(.A1(new_n697), .A2(new_n455), .A3(new_n699), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(G50gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g535(.A1(new_n637), .A2(new_n252), .A3(new_n702), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT107), .Z(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n687), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n458), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(G57gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  AOI21_X1  g541(.A(new_n459), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n687), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n675), .B2(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n546), .A2(new_n553), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g550(.A1(new_n739), .A2(new_n542), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n554), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n691), .A2(new_n693), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n253), .A2(new_n703), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT110), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n654), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n692), .B1(new_n686), .B2(new_n548), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(new_n757), .C1(KEYINPUT44), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n458), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n758), .B2(new_n756), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n429), .A2(new_n594), .A3(new_n654), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n759), .B2(new_n459), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n687), .A2(new_n688), .A3(new_n756), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT112), .A3(new_n761), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n346), .A2(new_n595), .A3(new_n654), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT111), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n767), .B(new_n779), .C1(new_n764), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n675), .B2(new_n759), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n677), .A2(G99gat), .A3(new_n702), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n764), .B2(new_n783), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n542), .A2(G106gat), .A3(new_n702), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n771), .A2(new_n773), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G106gat), .B1(new_n759), .B2(new_n542), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n762), .B2(new_n763), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(KEYINPUT113), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n786), .B2(new_n787), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n790), .A2(new_n787), .A3(new_n791), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1339gat));
  NAND4_X1  g597(.A1(new_n635), .A2(new_n253), .A3(new_n702), .A4(new_n636), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n241), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n233), .A2(new_n234), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n248), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT117), .A3(new_n654), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n641), .A2(new_n642), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n645), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n644), .A3(KEYINPUT54), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n812));
  OAI221_X1 g611(.A(new_n812), .B1(new_n643), .B2(new_n501), .C1(new_n641), .C2(new_n642), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n651), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n808), .B1(new_n814), .B2(new_n653), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n808), .A3(new_n653), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(new_n651), .A3(new_n813), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n816), .A2(new_n252), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n248), .A2(new_n654), .A3(new_n805), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n692), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n817), .A2(new_n820), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n815), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n688), .A3(new_n806), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n590), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT118), .B1(new_n801), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n799), .B(KEYINPUT114), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n703), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n455), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n346), .A2(new_n458), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n546), .A3(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(new_n354), .A3(new_n253), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n831), .A2(new_n836), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n543), .A2(new_n346), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n429), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n252), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n841), .A2(new_n846), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n840), .B2(new_n702), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n654), .A2(new_n368), .A3(new_n370), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n844), .B2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n840), .B2(new_n703), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n360), .A3(new_n590), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n836), .A3(new_n429), .ZN(new_n854));
  INV_X1    g653(.A(new_n843), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n688), .A2(new_n358), .ZN(new_n856));
  OR4_X1    g655(.A1(KEYINPUT119), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT119), .B1(new_n844), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n840), .B2(new_n692), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NAND4_X1  g663(.A1(new_n672), .A2(new_n455), .A3(new_n459), .A4(new_n673), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n253), .A2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n854), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT58), .B1(new_n868), .B2(KEYINPUT121), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n671), .A2(new_n839), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n831), .A2(new_n836), .A3(new_n455), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n829), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n252), .A2(new_n653), .A3(new_n814), .A4(new_n820), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n688), .B1(new_n878), .B2(new_n822), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n703), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n832), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n542), .A2(new_n875), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n873), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n386), .B1(new_n884), .B2(new_n252), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n870), .B1(new_n885), .B2(new_n868), .ZN(new_n886));
  INV_X1    g685(.A(new_n868), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n253), .B(new_n873), .C1(new_n876), .C2(new_n883), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n869), .B(new_n887), .C1(new_n888), .C2(new_n386), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n702), .B1(new_n873), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n799), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n799), .A2(new_n893), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n894), .A2(new_n880), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n875), .B1(new_n896), .B2(new_n542), .ZN(new_n897));
  INV_X1    g696(.A(new_n882), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n837), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n892), .B(new_n899), .C1(new_n891), .C2(new_n873), .ZN(new_n900));
  AND2_X1   g699(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n854), .A2(new_n865), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n702), .A2(G148gat), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n900), .A2(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n388), .B1(new_n884), .B2(new_n654), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(KEYINPUT59), .B2(new_n905), .ZN(G1345gat));
  INV_X1    g705(.A(G155gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n907), .A3(new_n590), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n884), .A2(new_n590), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n907), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n902), .B2(new_n688), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n688), .A2(G162gat), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n884), .B2(new_n912), .ZN(G1347gat));
  NOR4_X1   g712(.A1(new_n837), .A2(new_n429), .A3(new_n459), .A4(new_n543), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n273), .A3(new_n252), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n459), .A2(new_n429), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n677), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n838), .A2(new_n252), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(G169gat), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n919), .B2(G169gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n914), .B2(new_n654), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n842), .A2(new_n542), .A3(new_n918), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n654), .A2(new_n314), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n590), .A2(new_n277), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n914), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G183gat), .B1(new_n926), .B2(new_n703), .ZN(new_n933));
  XNOR2_X1  g732(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n914), .A2(new_n278), .A3(new_n688), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n838), .A2(new_n688), .A3(new_n918), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(G190gat), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n939), .B2(G190gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n674), .A2(new_n917), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n899), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(new_n253), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n672), .A2(new_n455), .A3(new_n346), .A4(new_n673), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n837), .A2(new_n429), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n252), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n948), .B1(new_n955), .B2(new_n947), .ZN(G1352gat));
  NOR2_X1   g755(.A1(new_n702), .A2(G204gat), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n951), .A2(new_n954), .A3(new_n952), .A4(new_n957), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n946), .B2(new_n702), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n899), .A2(new_n590), .A3(new_n945), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n953), .A2(new_n954), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n590), .A2(new_n261), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  OAI21_X1  g767(.A(G218gat), .B1(new_n946), .B2(new_n692), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n688), .A2(new_n262), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n966), .B2(new_n970), .ZN(G1355gat));
endmodule


