//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n204), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT93), .B(G29gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n203), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT94), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n203), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(KEYINPUT95), .B2(new_n207), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n207), .A2(KEYINPUT95), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT96), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT96), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(new_n213), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n211), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT97), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n230), .B(G8gat), .Z(new_n231));
  NOR2_X1   g030(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n231), .B1(new_n222), .B2(KEYINPUT17), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n233), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT98), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n234), .B(KEYINPUT13), .Z(new_n243));
  AND2_X1   g042(.A1(new_n222), .A2(new_n231), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(new_n232), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n221), .ZN(new_n246));
  INV_X1    g045(.A(new_n211), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n235), .A3(new_n231), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(new_n234), .A3(new_n233), .A4(new_n240), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n242), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G169gat), .B(G197gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n254), .A3(new_n261), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n266), .B1(KEYINPUT22), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n271), .B(new_n266), .C1(KEYINPUT22), .C2(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  AND2_X1   g081(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n283));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(KEYINPUT71), .B2(KEYINPUT26), .ZN(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  INV_X1    g085(.A(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT70), .B1(new_n288), .B2(KEYINPUT26), .ZN(new_n291));
  OAI221_X1 g090(.A(new_n282), .B1(new_n283), .B2(new_n285), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n281), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n284), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT65), .ZN(new_n306));
  OAI211_X1 g105(.A(KEYINPUT66), .B(new_n288), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT24), .B1(new_n293), .B2(KEYINPUT69), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(KEYINPUT69), .B2(new_n293), .ZN(new_n310));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n282), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n302), .B2(new_n307), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n293), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n293), .A2(KEYINPUT64), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT25), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n315), .B1(new_n324), .B2(KEYINPUT67), .ZN(new_n325));
  INV_X1    g124(.A(new_n316), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n301), .A2(new_n300), .A3(new_n284), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n305), .A2(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT66), .B1(new_n330), .B2(new_n288), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n323), .B(new_n326), .C1(new_n327), .C2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT67), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n294), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n276), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT67), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n334), .A3(new_n315), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n275), .B1(new_n342), .B2(new_n294), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n273), .B(new_n274), .C1(new_n338), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n276), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n273), .A2(new_n274), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n342), .B2(new_n294), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n276), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT37), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT89), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT38), .ZN(new_n355));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n344), .A2(new_n348), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT37), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n354), .B2(new_n360), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  INV_X1    g163(.A(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G113gat), .A2(G120gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n371), .A3(new_n367), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n372), .B(new_n363), .C1(new_n368), .C2(new_n369), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT77), .B1(new_n378), .B2(G141gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380));
  INV_X1    g179(.A(G141gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(G148gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(G141gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT78), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n379), .A2(new_n382), .A3(new_n386), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n385), .A2(new_n387), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n381), .A2(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n383), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n390), .ZN(new_n395));
  INV_X1    g194(.A(new_n388), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n377), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n387), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n388), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n376), .A3(new_n398), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT79), .B(KEYINPUT5), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n400), .B2(new_n404), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n403), .A2(new_n412), .A3(new_n398), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(new_n392), .B2(new_n399), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n377), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n392), .A2(new_n399), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n415), .A2(new_n417), .A3(new_n406), .A4(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n407), .A2(new_n411), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT80), .ZN(new_n422));
  INV_X1    g221(.A(new_n420), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n420), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n421), .B(new_n430), .C1(new_n424), .C2(new_n425), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n344), .A2(new_n348), .A3(new_n358), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT76), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT76), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n344), .A2(new_n348), .A3(new_n439), .A4(new_n358), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n361), .A2(new_n362), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n443), .B(KEYINPUT83), .Z(new_n444));
  AOI21_X1  g243(.A(new_n346), .B1(new_n413), .B2(new_n337), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT3), .B1(new_n346), .B2(new_n337), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n418), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n444), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT29), .B1(new_n418), .B2(new_n412), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n449), .A2(new_n346), .B1(new_n418), .B2(new_n446), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n448), .A2(KEYINPUT84), .B1(new_n450), .B2(new_n443), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(new_n444), .ZN(new_n453));
  OAI21_X1  g252(.A(G22gat), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n452), .A3(new_n444), .ZN(new_n456));
  INV_X1    g255(.A(G22gat), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n445), .A2(new_n447), .A3(new_n443), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n454), .A2(new_n465), .A3(new_n459), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n454), .A2(new_n459), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n462), .B(KEYINPUT82), .Z(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(KEYINPUT85), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT85), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n438), .A2(new_n474), .A3(new_n440), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n358), .B1(new_n344), .B2(new_n348), .ZN(new_n476));
  INV_X1    g275(.A(new_n437), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(KEYINPUT30), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n415), .A2(new_n417), .A3(new_n419), .ZN(new_n481));
  INV_X1    g280(.A(new_n406), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n480), .B1(new_n405), .B2(new_n406), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n485), .A2(new_n491), .A3(KEYINPUT40), .A4(new_n430), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n432), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n485), .A2(new_n491), .A3(new_n430), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n473), .B1(new_n479), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT90), .B1(new_n442), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n468), .A2(new_n469), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n504), .A2(new_n470), .B1(new_n464), .B2(new_n466), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n432), .A2(new_n492), .ZN(new_n506));
  INV_X1    g305(.A(new_n498), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n475), .A2(new_n478), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n354), .A2(new_n360), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n435), .A2(new_n436), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n438), .A2(new_n440), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n434), .A2(new_n433), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n434), .A2(KEYINPUT81), .A3(new_n433), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n432), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n436), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n473), .B1(new_n526), .B2(new_n479), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n529));
  NAND2_X1  g328(.A1(G227gat), .A2(G233gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n294), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n339), .A2(new_n340), .B1(new_n314), .B2(new_n308), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n376), .B(new_n531), .C1(new_n532), .C2(new_n334), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n377), .B1(new_n342), .B2(new_n294), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT75), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n336), .A2(new_n376), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n342), .A2(new_n377), .A3(new_n294), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT75), .A3(new_n529), .A4(new_n530), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT34), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n537), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n530), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n538), .A2(new_n545), .A3(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G43gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT74), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G99gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n546), .B2(KEYINPUT32), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n546), .B(KEYINPUT32), .C1(new_n547), .C2(new_n555), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n544), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n545), .B1(new_n538), .B2(new_n539), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT75), .B1(new_n560), .B2(new_n529), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n529), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n557), .A2(new_n558), .B1(new_n563), .B2(new_n541), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT36), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n558), .ZN(new_n566));
  INV_X1    g365(.A(new_n544), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n544), .A2(new_n557), .A3(new_n558), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n520), .A2(new_n528), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n559), .A2(new_n564), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n526), .A3(new_n473), .A4(new_n479), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n514), .A2(new_n510), .A3(KEYINPUT35), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n570), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n505), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n575), .A2(KEYINPUT35), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n265), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n526), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n585), .A2(new_n591), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n231), .B1(new_n584), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT100), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n584), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT99), .Z(new_n599));
  XOR2_X1   g398(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G183gat), .B(G211gat), .Z(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n609), .A3(new_n603), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n615), .B(new_n617), .Z(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT103), .Z(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(G85gat), .ZN(new_n622));
  INV_X1    g421(.A(G92gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(KEYINPUT8), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(KEYINPUT102), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT7), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n621), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n621), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n624), .A2(new_n632), .A3(new_n625), .A4(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n250), .A2(new_n235), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n248), .A2(new_n636), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n620), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n618), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n620), .A3(new_n637), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n638), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n644), .A2(new_n639), .A3(new_n641), .A4(new_n618), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n634), .B(new_n595), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT106), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n634), .A2(new_n595), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT105), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n650), .A2(KEYINPUT10), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n656), .A2(KEYINPUT105), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n651), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n649), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n649), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT107), .B(new_n664), .C1(new_n654), .C2(new_n660), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n613), .A2(new_n646), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n583), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(G1gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n581), .A2(new_n510), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n668), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G8gat), .B1(new_n673), .B2(new_n668), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n672), .A2(KEYINPUT109), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n676), .A2(new_n677), .B1(new_n674), .B2(new_n681), .ZN(G1325gat));
  INV_X1    g481(.A(new_n668), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n565), .A2(KEYINPUT110), .A3(new_n571), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT110), .B1(new_n565), .B2(new_n571), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n581), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n581), .A2(new_n574), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n668), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(G1326gat));
  INV_X1    g491(.A(new_n265), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n528), .A2(new_n572), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n501), .B2(new_n519), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n693), .B(new_n505), .C1(new_n695), .C2(new_n579), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n668), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n613), .A2(new_n646), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n667), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n209), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n583), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n581), .A2(KEYINPUT45), .A3(new_n582), .A4(new_n703), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n684), .A2(new_n685), .A3(new_n527), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n579), .B1(new_n520), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n646), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n646), .A2(new_n707), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n695), .B2(new_n579), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n666), .B(KEYINPUT111), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n613), .A3(new_n265), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n582), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n209), .B1(new_n717), .B2(new_n718), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n705), .B(new_n706), .C1(new_n719), .C2(new_n720), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n713), .A2(new_n510), .A3(new_n716), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G36gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n702), .A2(G36gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT46), .B1(new_n673), .B2(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n673), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(G1329gat));
  OR2_X1    g527(.A1(new_n702), .A2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n690), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n710), .A2(new_n687), .A3(new_n712), .A4(new_n716), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(G43gat), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n710), .A2(new_n505), .A3(new_n712), .A4(new_n716), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(new_n735), .A3(G50gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n734), .B2(G50gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n702), .A2(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n696), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT48), .B1(new_n696), .B2(new_n739), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n734), .B2(G50gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT114), .B(new_n742), .C1(new_n734), .C2(G50gat), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n741), .A2(KEYINPUT48), .B1(new_n745), .B2(new_n746), .ZN(G1331gat));
  NOR2_X1   g546(.A1(new_n709), .A2(new_n693), .ZN(new_n748));
  INV_X1    g547(.A(new_n613), .ZN(new_n749));
  INV_X1    g548(.A(new_n646), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n749), .A2(new_n750), .A3(new_n714), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n526), .B(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT116), .B(G57gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n510), .A3(new_n751), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  XNOR2_X1  g561(.A(new_n577), .B(KEYINPUT117), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n748), .A2(new_n751), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n687), .A2(G71gat), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n764), .A2(G71gat), .B1(new_n752), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n473), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n588), .ZN(G1335gat));
  NOR3_X1   g568(.A1(new_n693), .A2(new_n613), .A3(new_n667), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n713), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n526), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT51), .B1(new_n748), .B2(new_n701), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n701), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n582), .A2(new_n622), .A3(new_n666), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NOR3_X1   g578(.A1(new_n714), .A2(G92gat), .A3(new_n479), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n710), .A2(new_n510), .A3(new_n712), .A4(new_n770), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n780), .B(KEYINPUT118), .Z(new_n786));
  AOI22_X1  g585(.A1(new_n776), .A2(new_n786), .B1(G92gat), .B2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n771), .B2(new_n686), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n577), .A2(G99gat), .A3(new_n667), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n777), .B2(new_n790), .ZN(G1338gat));
  NOR2_X1   g590(.A1(new_n714), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n775), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n505), .B(new_n792), .C1(new_n793), .C2(new_n773), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n710), .A2(new_n505), .A3(new_n712), .A4(new_n770), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1339gat));
  INV_X1    g600(.A(new_n578), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n242), .A2(new_n252), .A3(new_n245), .A4(new_n261), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n234), .B1(new_n251), .B2(new_n233), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n244), .A2(new_n232), .A3(new_n243), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n260), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n666), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n660), .A2(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n649), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n652), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .A3(new_n660), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n809), .B2(new_n812), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n661), .A2(new_n664), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n646), .B(new_n807), .C1(new_n265), .C2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n815), .A2(new_n818), .A3(new_n806), .A4(new_n803), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n613), .B1(new_n821), .B2(new_n750), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n683), .A2(new_n265), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n802), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n526), .A2(new_n510), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n364), .A3(new_n265), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n829), .A2(KEYINPUT121), .A3(new_n754), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT121), .B1(new_n829), .B2(new_n754), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n693), .B(new_n479), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n835), .B2(new_n364), .ZN(G1340gat));
  NOR3_X1   g635(.A1(new_n831), .A2(new_n365), .A3(new_n714), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n666), .B(new_n479), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n365), .ZN(G1341gat));
  NOR2_X1   g638(.A1(new_n749), .A2(G127gat), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n479), .B(new_n840), .C1(new_n833), .C2(new_n834), .ZN(new_n841));
  OAI21_X1  g640(.A(G127gat), .B1(new_n831), .B2(new_n749), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NOR2_X1   g642(.A1(new_n646), .A2(new_n510), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT122), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(G134gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n833), .B2(new_n834), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n831), .B2(new_n646), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  AOI21_X1  g650(.A(new_n473), .B1(new_n826), .B2(new_n828), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(new_n479), .A3(new_n686), .A4(new_n754), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n381), .B1(new_n853), .B2(new_n265), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n686), .A2(new_n830), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n825), .A2(new_n505), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n265), .A2(new_n381), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n854), .B(KEYINPUT58), .C1(new_n861), .C2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1344gat));
  AND3_X1   g667(.A1(new_n823), .A2(new_n827), .A3(new_n824), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n827), .B1(new_n823), .B2(new_n824), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT57), .B(new_n505), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n859), .A2(new_n855), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n858), .A2(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n858), .A2(KEYINPUT123), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n666), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT59), .B(G148gat), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n826), .A2(new_n828), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n505), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n687), .A3(new_n755), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n880), .A2(new_n378), .A3(new_n666), .A4(new_n479), .ZN(new_n881));
  INV_X1    g680(.A(new_n861), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n378), .B1(new_n882), .B2(new_n666), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n877), .B(new_n881), .C1(new_n883), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n861), .B2(new_n749), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n749), .A2(G155gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n853), .B2(new_n886), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n861), .B2(new_n646), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n845), .A2(G162gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n754), .A2(new_n479), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n473), .A3(new_n763), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n286), .A3(new_n265), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n582), .A2(new_n479), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n829), .A2(new_n693), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n286), .B2(new_n897), .ZN(G1348gat));
  OAI21_X1  g697(.A(G176gat), .B1(new_n894), .B2(new_n714), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n829), .A2(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n666), .A2(new_n287), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g702(.A(G183gat), .B1(new_n894), .B2(new_n749), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n613), .A2(new_n277), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n878), .A2(new_n750), .A3(new_n893), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G190gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n911), .A3(G190gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n912), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n829), .A2(new_n278), .A3(new_n750), .A4(new_n896), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT125), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n879), .A2(new_n687), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n693), .A3(new_n896), .ZN(new_n921));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n892), .A2(new_n686), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n871), .B2(new_n872), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n265), .A2(new_n922), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n921), .A2(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n667), .A2(G204gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n920), .A2(new_n896), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT62), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT62), .ZN(new_n930));
  INV_X1    g729(.A(G204gat), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n924), .A2(new_n715), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(G1353gat));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n924), .A2(new_n613), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n267), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n920), .A2(new_n267), .A3(new_n613), .A4(new_n896), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n267), .B1(new_n924), .B2(new_n613), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(new_n939), .B2(KEYINPUT63), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n935), .B(new_n267), .C1(new_n924), .C2(new_n613), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n937), .B(new_n938), .C1(new_n940), .C2(new_n941), .ZN(G1354gat));
  AND2_X1   g741(.A1(new_n924), .A2(new_n750), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n896), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n750), .A2(new_n268), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n943), .A2(new_n268), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


