

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U550 ( .A1(n707), .A2(n518), .ZN(n708) );
  OR2_X1 U551 ( .A1(n588), .A2(n775), .ZN(n589) );
  AND2_X2 U552 ( .A1(n523), .A2(G2104), .ZN(n580) );
  NAND2_X1 U553 ( .A1(n591), .A2(n732), .ZN(n654) );
  INV_X2 U554 ( .A(G2105), .ZN(n523) );
  AND2_X1 U555 ( .A1(n709), .A2(n708), .ZN(n710) );
  BUF_X1 U556 ( .A(n715), .Z(n716) );
  XNOR2_X2 U557 ( .A(n590), .B(KEYINPUT92), .ZN(n731) );
  AND2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n890) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(n519), .Z(n715) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  BUF_X1 U561 ( .A(n654), .Z(n667) );
  NOR2_X1 U562 ( .A1(n706), .A2(n688), .ZN(n689) );
  NOR2_X1 U563 ( .A1(n562), .A2(G651), .ZN(n529) );
  INV_X1 U564 ( .A(KEYINPUT23), .ZN(n581) );
  AND2_X1 U565 ( .A1(n526), .A2(n515), .ZN(G164) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n523), .ZN(n585) );
  AND2_X1 U567 ( .A1(n525), .A2(n524), .ZN(n515) );
  XOR2_X1 U568 ( .A(n645), .B(KEYINPUT28), .Z(n516) );
  AND2_X1 U569 ( .A1(n934), .A2(n760), .ZN(n517) );
  OR2_X1 U570 ( .A1(n706), .A2(n705), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n679), .A2(n656), .ZN(n658) );
  INV_X1 U572 ( .A(KEYINPUT29), .ZN(n647) );
  INV_X1 U573 ( .A(n919), .ZN(n688) );
  INV_X1 U574 ( .A(KEYINPUT32), .ZN(n675) );
  AND2_X1 U575 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U576 ( .A(n621), .B(KEYINPUT76), .ZN(n622) );
  NOR2_X1 U577 ( .A1(n744), .A2(n517), .ZN(n745) );
  XNOR2_X1 U578 ( .A(n623), .B(n622), .ZN(n636) );
  BUF_X1 U579 ( .A(n636), .Z(n937) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n562) );
  XNOR2_X1 U581 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U582 ( .A(n522), .B(KEYINPUT91), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT67), .B(n540), .Z(G171) );
  NAND2_X1 U584 ( .A1(G102), .A2(n580), .ZN(n521) );
  NAND2_X1 U585 ( .A1(G138), .A2(n715), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U587 ( .A1(G114), .A2(n890), .ZN(n525) );
  NAND2_X1 U588 ( .A1(G126), .A2(n585), .ZN(n524) );
  INV_X1 U589 ( .A(G651), .ZN(n533) );
  NOR2_X1 U590 ( .A1(G543), .A2(n533), .ZN(n527) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n527), .Z(n790) );
  NAND2_X1 U592 ( .A1(G64), .A2(n790), .ZN(n531) );
  INV_X1 U593 ( .A(KEYINPUT65), .ZN(n528) );
  XNOR2_X2 U594 ( .A(n529), .B(n528), .ZN(n791) );
  NAND2_X1 U595 ( .A1(G52), .A2(n791), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n539) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n794) );
  NAND2_X1 U598 ( .A1(n794), .A2(G90), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT66), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n562), .A2(n533), .ZN(n534) );
  NAND2_X1 U601 ( .A1(G77), .A2(n534), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n537), .Z(n538) );
  NOR2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U605 ( .A1(G63), .A2(n790), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G51), .A2(n791), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n543), .Z(n551) );
  NAND2_X1 U609 ( .A1(G76), .A2(n534), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT77), .B(KEYINPUT4), .Z(n545) );
  NAND2_X1 U611 ( .A1(G89), .A2(n794), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT5), .ZN(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT78), .B(n549), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n552), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G75), .A2(n534), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G88), .A2(n794), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G62), .A2(n790), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G50), .A2(n791), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(G166) );
  INV_X1 U626 ( .A(G166), .ZN(G303) );
  NAND2_X1 U627 ( .A1(G49), .A2(n791), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U630 ( .A1(n790), .A2(n561), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n562), .A2(G87), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(G288) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n566) );
  NAND2_X1 U634 ( .A1(G73), .A2(n534), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n566), .B(n565), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G61), .A2(n790), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G86), .A2(n794), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n791), .A2(G48), .ZN(n569) );
  XOR2_X1 U640 ( .A(KEYINPUT84), .B(n569), .Z(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(G305) );
  AND2_X1 U643 ( .A1(n790), .A2(G60), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G72), .A2(n534), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G85), .A2(n794), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n791), .A2(G47), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(G290) );
  NAND2_X1 U650 ( .A1(n715), .A2(G137), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G101), .A2(n580), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n776) );
  INV_X1 U653 ( .A(G40), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G113), .A2(n890), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G125), .A2(n585), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n775) );
  OR2_X2 U657 ( .A1(n776), .A2(n589), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n731), .B(KEYINPUT97), .ZN(n591) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n732) );
  INV_X2 U660 ( .A(n654), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n593), .A2(G2072), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT27), .ZN(n595) );
  INV_X1 U663 ( .A(G1956), .ZN(n945) );
  NOR2_X1 U664 ( .A1(n945), .A2(n593), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n644) );
  NAND2_X1 U666 ( .A1(G91), .A2(n794), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G53), .A2(n791), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G65), .A2(n790), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G78), .A2(n534), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT68), .ZN(n931) );
  NAND2_X1 U674 ( .A1(n644), .A2(n931), .ZN(n643) );
  NAND2_X1 U675 ( .A1(n790), .A2(G56), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT14), .B(n603), .Z(n611) );
  NAND2_X1 U677 ( .A1(G68), .A2(n534), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT71), .B(KEYINPUT12), .Z(n605) );
  NAND2_X1 U679 ( .A1(G81), .A2(n794), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT13), .ZN(n609) );
  XOR2_X1 U683 ( .A(KEYINPUT72), .B(n609), .Z(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n791), .A2(G43), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n932) );
  NAND2_X1 U687 ( .A1(G54), .A2(n791), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G79), .A2(n534), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT75), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G66), .A2(n790), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G92), .A2(n794), .ZN(n617) );
  AND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n623) );
  INV_X1 U695 ( .A(KEYINPUT15), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n636), .A2(G1348), .ZN(n626) );
  INV_X1 U697 ( .A(G1341), .ZN(n624) );
  AND2_X1 U698 ( .A1(n624), .A2(KEYINPUT26), .ZN(n625) );
  AND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U700 ( .A1(n627), .A2(n593), .ZN(n628) );
  OR2_X1 U701 ( .A1(n932), .A2(n628), .ZN(n635) );
  NAND2_X1 U702 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n636), .A2(G2067), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n593), .A2(n631), .ZN(n633) );
  OR2_X1 U706 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n641) );
  NAND2_X1 U709 ( .A1(G1348), .A2(n667), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G2067), .A2(n593), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U712 ( .A1(n937), .A2(n639), .ZN(n640) );
  NOR2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n644), .A2(n931), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n516), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n653) );
  XOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .Z(n1000) );
  NAND2_X1 U719 ( .A1(n593), .A2(n1000), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G1961), .A2(n667), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT100), .B(n651), .Z(n660) );
  NAND2_X1 U723 ( .A1(n660), .A2(G171), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n665) );
  NAND2_X1 U725 ( .A1(G8), .A2(n654), .ZN(n706) );
  NOR2_X1 U726 ( .A1(G1966), .A2(n706), .ZN(n679) );
  NOR2_X2 U727 ( .A1(n654), .A2(G2084), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT99), .ZN(n677) );
  NAND2_X1 U729 ( .A1(G8), .A2(n677), .ZN(n656) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(KEYINPUT101), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U732 ( .A1(G168), .A2(n659), .ZN(n662) );
  NOR2_X1 U733 ( .A1(G171), .A2(n660), .ZN(n661) );
  NOR2_X2 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT31), .B(n663), .Z(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT102), .ZN(n680) );
  NAND2_X1 U738 ( .A1(n680), .A2(G286), .ZN(n674) );
  INV_X1 U739 ( .A(G8), .ZN(n672) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n706), .ZN(n669) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G303), .ZN(n671) );
  OR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n676), .B(n675), .ZN(n685) );
  INV_X1 U747 ( .A(n677), .ZN(n678) );
  NAND2_X1 U748 ( .A1(G8), .A2(n678), .ZN(n683) );
  INV_X1 U749 ( .A(n679), .ZN(n681) );
  AND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n699) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n694) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n694), .A2(n686), .ZN(n920) );
  XOR2_X1 U756 ( .A(n920), .B(KEYINPUT103), .Z(n687) );
  NAND2_X1 U757 ( .A1(n699), .A2(n687), .ZN(n690) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n919) );
  XNOR2_X1 U759 ( .A(n691), .B(KEYINPUT64), .ZN(n692) );
  NOR2_X1 U760 ( .A1(KEYINPUT33), .A2(n692), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n693), .B(KEYINPUT104), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n694), .A2(KEYINPUT33), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n706), .A2(n695), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n926) );
  NAND2_X1 U766 ( .A1(n698), .A2(n926), .ZN(n709) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n700) );
  NAND2_X1 U768 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n699), .A2(n701), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n702), .A2(n706), .ZN(n707) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U772 ( .A(n703), .B(KEYINPUT98), .Z(n704) );
  XNOR2_X1 U773 ( .A(KEYINPUT24), .B(n704), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT105), .ZN(n746) );
  NAND2_X1 U775 ( .A1(n585), .A2(G119), .ZN(n711) );
  XOR2_X1 U776 ( .A(KEYINPUT93), .B(n711), .Z(n713) );
  NAND2_X1 U777 ( .A1(n890), .A2(G107), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U779 ( .A(KEYINPUT94), .B(n714), .Z(n718) );
  NAND2_X1 U780 ( .A1(n716), .A2(G131), .ZN(n717) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U782 ( .A1(G95), .A2(n580), .ZN(n719) );
  XNOR2_X1 U783 ( .A(KEYINPUT95), .B(n719), .ZN(n720) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n882) );
  INV_X1 U785 ( .A(G1991), .ZN(n749) );
  NOR2_X1 U786 ( .A1(n882), .A2(n749), .ZN(n730) );
  INV_X1 U787 ( .A(G1996), .ZN(n999) );
  NAND2_X1 U788 ( .A1(n580), .A2(G105), .ZN(n722) );
  XNOR2_X1 U789 ( .A(n722), .B(KEYINPUT38), .ZN(n724) );
  NAND2_X1 U790 ( .A1(G141), .A2(n716), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U792 ( .A1(G117), .A2(n890), .ZN(n726) );
  NAND2_X1 U793 ( .A1(G129), .A2(n585), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U795 ( .A1(n728), .A2(n727), .ZN(n877) );
  NOR2_X1 U796 ( .A1(n999), .A2(n877), .ZN(n729) );
  NOR2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n979) );
  NOR2_X1 U798 ( .A1(n731), .A2(n732), .ZN(n760) );
  XOR2_X1 U799 ( .A(n760), .B(KEYINPUT96), .Z(n733) );
  NOR2_X1 U800 ( .A1(n979), .A2(n733), .ZN(n752) );
  INV_X1 U801 ( .A(n752), .ZN(n743) );
  NAND2_X1 U802 ( .A1(G116), .A2(n890), .ZN(n735) );
  NAND2_X1 U803 ( .A1(G128), .A2(n585), .ZN(n734) );
  NAND2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U805 ( .A(n736), .B(KEYINPUT35), .ZN(n741) );
  NAND2_X1 U806 ( .A1(G104), .A2(n580), .ZN(n738) );
  NAND2_X1 U807 ( .A1(G140), .A2(n716), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U809 ( .A(KEYINPUT34), .B(n739), .Z(n740) );
  NAND2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U811 ( .A(n742), .B(KEYINPUT36), .Z(n878) );
  XNOR2_X1 U812 ( .A(KEYINPUT37), .B(G2067), .ZN(n747) );
  NOR2_X1 U813 ( .A1(n878), .A2(n747), .ZN(n977) );
  NAND2_X1 U814 ( .A1(n760), .A2(n977), .ZN(n758) );
  NAND2_X1 U815 ( .A1(n743), .A2(n758), .ZN(n744) );
  XNOR2_X1 U816 ( .A(G1986), .B(G290), .ZN(n934) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n763) );
  AND2_X1 U818 ( .A1(n878), .A2(n747), .ZN(n748) );
  XOR2_X1 U819 ( .A(KEYINPUT108), .B(n748), .Z(n984) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n750) );
  AND2_X1 U821 ( .A1(n749), .A2(n882), .ZN(n981) );
  NOR2_X1 U822 ( .A1(n750), .A2(n981), .ZN(n751) );
  NOR2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n754) );
  AND2_X1 U824 ( .A1(n877), .A2(n999), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT106), .ZN(n986) );
  NOR2_X1 U826 ( .A1(n754), .A2(n986), .ZN(n756) );
  XOR2_X1 U827 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n755) );
  XNOR2_X1 U828 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n984), .A2(n759), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U832 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U833 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U835 ( .A1(G135), .A2(n716), .ZN(n766) );
  NAND2_X1 U836 ( .A1(G111), .A2(n890), .ZN(n765) );
  NAND2_X1 U837 ( .A1(n766), .A2(n765), .ZN(n771) );
  XOR2_X1 U838 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n768) );
  NAND2_X1 U839 ( .A1(G123), .A2(n585), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U841 ( .A(KEYINPUT80), .B(n769), .Z(n770) );
  NOR2_X1 U842 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U843 ( .A1(n580), .A2(G99), .ZN(n772) );
  NAND2_X1 U844 ( .A1(n773), .A2(n772), .ZN(n974) );
  XNOR2_X1 U845 ( .A(G2096), .B(n974), .ZN(n774) );
  OR2_X1 U846 ( .A1(G2100), .A2(n774), .ZN(G156) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  INV_X1 U849 ( .A(G69), .ZN(G235) );
  INV_X1 U850 ( .A(G108), .ZN(G238) );
  INV_X1 U851 ( .A(G120), .ZN(G236) );
  NOR2_X1 U852 ( .A1(n776), .A2(n775), .ZN(G160) );
  NAND2_X1 U853 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U854 ( .A(n777), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U855 ( .A(G223), .ZN(n833) );
  NAND2_X1 U856 ( .A1(n833), .A2(G567), .ZN(n778) );
  XOR2_X1 U857 ( .A(KEYINPUT11), .B(n778), .Z(G234) );
  INV_X1 U858 ( .A(G860), .ZN(n801) );
  OR2_X1 U859 ( .A1(n932), .A2(n801), .ZN(G153) );
  XNOR2_X1 U860 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n779) );
  XNOR2_X1 U862 ( .A(n779), .B(KEYINPUT74), .ZN(n781) );
  INV_X1 U863 ( .A(G868), .ZN(n813) );
  NAND2_X1 U864 ( .A1(n937), .A2(n813), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G284) );
  XNOR2_X1 U866 ( .A(KEYINPUT69), .B(n931), .ZN(G299) );
  NOR2_X1 U867 ( .A1(G286), .A2(n813), .ZN(n782) );
  XOR2_X1 U868 ( .A(KEYINPUT79), .B(n782), .Z(n784) );
  NOR2_X1 U869 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U871 ( .A1(n801), .A2(G559), .ZN(n785) );
  INV_X1 U872 ( .A(n937), .ZN(n799) );
  NAND2_X1 U873 ( .A1(n785), .A2(n799), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U875 ( .A1(G868), .A2(n932), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n799), .A2(G868), .ZN(n787) );
  NOR2_X1 U877 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U879 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U880 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G80), .A2(n534), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G93), .A2(n794), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n812) );
  XOR2_X1 U886 ( .A(n812), .B(KEYINPUT82), .Z(n803) );
  NAND2_X1 U887 ( .A1(n799), .A2(G559), .ZN(n800) );
  XOR2_X1 U888 ( .A(n932), .B(n800), .Z(n810) );
  NAND2_X1 U889 ( .A1(n810), .A2(n801), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n803), .B(n802), .ZN(G145) );
  XNOR2_X1 U891 ( .A(G166), .B(G290), .ZN(n809) );
  XNOR2_X1 U892 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n805) );
  XNOR2_X1 U893 ( .A(G288), .B(G299), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n812), .B(n806), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n807), .B(G305), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n898) );
  XNOR2_X1 U898 ( .A(n810), .B(n898), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n811), .A2(G868), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT86), .B(n816), .Z(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n817), .Z(n818) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XOR2_X1 U908 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U909 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U910 ( .A1(G236), .A2(G238), .ZN(n822) );
  NOR2_X1 U911 ( .A1(G235), .A2(G237), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U913 ( .A(KEYINPUT88), .B(n823), .ZN(n838) );
  NAND2_X1 U914 ( .A1(G567), .A2(n838), .ZN(n829) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n824), .Z(n825) );
  NOR2_X1 U917 ( .A1(G218), .A2(n825), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G96), .A2(n826), .ZN(n837) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n837), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT87), .B(n827), .Z(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n839) );
  NAND2_X1 U922 ( .A1(G661), .A2(G483), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT89), .B(n830), .Z(n831) );
  NOR2_X1 U924 ( .A1(n839), .A2(n831), .ZN(n836) );
  NAND2_X1 U925 ( .A1(G36), .A2(n836), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n832), .B(KEYINPUT90), .ZN(G176) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U932 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  INV_X1 U936 ( .A(n839), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2678), .B(G2084), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2078), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n842), .B(G2100), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2072), .B(G2090), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(G2096), .B(KEYINPUT111), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1981), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1961), .B(G1956), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n851), .B(G2474), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1966), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1971), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n585), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G100), .A2(n580), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n859), .B(KEYINPUT112), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G136), .A2(n716), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G112), .A2(n890), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n875) );
  NAND2_X1 U967 ( .A1(G103), .A2(n580), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G139), .A2(n716), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G115), .A2(n890), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G127), .A2(n585), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(n871), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n970) );
  XNOR2_X1 U976 ( .A(n970), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(n876), .B(G162), .Z(n880) );
  XOR2_X1 U979 ( .A(n878), .B(n877), .Z(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n974), .B(n881), .ZN(n884) );
  XNOR2_X1 U982 ( .A(G160), .B(n882), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G106), .A2(n580), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G142), .A2(n716), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n887), .B(KEYINPUT45), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G130), .A2(n585), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G118), .A2(n890), .ZN(n891) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n891), .ZN(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(G164), .B(n894), .Z(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n932), .B(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(G171), .B(n937), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(G286), .B(n901), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2451), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G2446), .B(G2427), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n911) );
  XOR2_X1 U1004 ( .A(G2438), .B(KEYINPUT109), .Z(n906) );
  XNOR2_X1 U1005 ( .A(G2443), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1007 ( .A(n907), .B(G2435), .Z(n909) );
  XNOR2_X1 U1008 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .ZN(n943) );
  NAND2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n922) );
  AND2_X1 U1023 ( .A1(G303), .A2(G1971), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1025 ( .A(KEYINPUT123), .B(n923), .Z(n925) );
  XNOR2_X1 U1026 ( .A(G171), .B(G1961), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1030 ( .A(KEYINPUT57), .B(n928), .Z(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G1956), .B(n931), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G1341), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1348), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT124), .B(n944), .ZN(n1026) );
  XNOR2_X1 U1041 ( .A(G20), .B(n945), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G6), .B(G1981), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1046 ( .A(KEYINPUT59), .B(G1348), .Z(n950) );
  XNOR2_X1 U1047 ( .A(G4), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n953), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(G1986), .B(G24), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1057 ( .A(G1971), .B(KEYINPUT126), .Z(n960) );
  XNOR2_X1 U1058 ( .A(G22), .B(n960), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n966), .B(KEYINPUT61), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT125), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n969), .ZN(n1024) );
  INV_X1 U1066 ( .A(KEYINPUT55), .ZN(n996) );
  XOR2_X1 U1067 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(KEYINPUT50), .B(n973), .ZN(n993) );
  XNOR2_X1 U1071 ( .A(G160), .B(G2084), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT116), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G2090), .B(G162), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT117), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1085 ( .A(KEYINPUT52), .B(n994), .Z(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1088 ( .A(G2084), .B(G34), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT54), .ZN(n1017) );
  XNOR2_X1 U1090 ( .A(G2090), .B(G35), .ZN(n1014) );
  XNOR2_X1 U1091 ( .A(G32), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n1000), .B(G27), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G2072), .B(G33), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT119), .B(G2067), .Z(n1005) );
  XNOR2_X1 U1097 ( .A(G26), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(KEYINPUT120), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(G28), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(G25), .B(G1991), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(KEYINPUT121), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT55), .B(n1018), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(KEYINPUT122), .B(n1020), .Z(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(n1028), .B(n1027), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

