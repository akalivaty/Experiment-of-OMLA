//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g0039(.A1(G68), .A2(G77), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n203), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G351));
  AOI21_X1  g0045(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n206), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G226), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n256), .B(new_n206), .C1(new_n261), .C2(G45), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G222), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G223), .A3(G1698), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(new_n202), .C2(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n246), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g0072(.A(KEYINPUT70), .B(G179), .Z(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n277), .A2(new_n215), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n207), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n276), .B1(new_n280), .B2(G50), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g0084(.A(G58), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n285), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n284), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n207), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G150), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n294), .A2(new_n296), .B1(new_n297), .B2(new_n207), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n277), .A2(new_n215), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n282), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n274), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT66), .B(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n251), .A2(G244), .B1(new_n306), .B2(new_n256), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  OAI211_X1 g0109(.A(G232), .B(new_n265), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(G238), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n311));
  OR2_X1    g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G107), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n246), .ZN(new_n316));
  AOI21_X1  g0116(.A(G169), .B1(new_n307), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n275), .A2(G77), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n279), .B2(new_n202), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G20), .A2(G77), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n321), .B1(new_n283), .B2(new_n296), .C1(new_n291), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n301), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT71), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n315), .A2(new_n246), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n254), .A2(new_n255), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n257), .A2(new_n305), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT67), .B1(new_n328), .B2(new_n206), .ZN(new_n329));
  INV_X1    g0129(.A(new_n250), .ZN(new_n330));
  OAI211_X1 g0130(.A(G244), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n262), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n271), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n320), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(new_n301), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n273), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n307), .A2(new_n339), .A3(new_n316), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n325), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n307), .A2(new_n316), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n336), .B1(G200), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n342), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n303), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n228), .A2(G1698), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G226), .B2(G1698), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n308), .A2(new_n309), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n246), .B1(new_n306), .B2(new_n256), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n251), .A2(G238), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(G190), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n202), .B2(new_n291), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n360), .A2(KEYINPUT11), .A3(new_n301), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT12), .ZN(new_n362));
  INV_X1    g0162(.A(new_n275), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n201), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n275), .A2(KEYINPUT12), .A3(G68), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n279), .A2(new_n201), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT11), .B1(new_n360), .B2(new_n301), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n355), .B2(new_n357), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n357), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n355), .A2(G179), .A3(new_n357), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n377), .A3(G169), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n368), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n284), .A2(new_n289), .A3(new_n286), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n289), .B1(new_n284), .B2(new_n286), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n363), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n288), .A2(new_n290), .A3(new_n280), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n350), .B2(new_n207), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n308), .A2(new_n309), .A3(new_n388), .A4(G20), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n285), .A2(new_n201), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n295), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n278), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n386), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G226), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G223), .B2(G1698), .ZN(new_n404));
  INV_X1    g0204(.A(G33), .ZN(new_n405));
  INV_X1    g0205(.A(G87), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n404), .A2(new_n350), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n246), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n251), .A2(G232), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n262), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n271), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n273), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT18), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n410), .A2(new_n271), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n410), .A2(new_n273), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n384), .A2(new_n385), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n388), .B1(new_n264), .B2(G20), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n350), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n201), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n398), .B1(new_n420), .B2(new_n395), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n400), .A3(new_n301), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n413), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n402), .B2(G1698), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n264), .B1(G33), .B2(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n262), .B1(new_n429), .B2(new_n327), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n251), .A2(G232), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n370), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n408), .A2(new_n409), .A3(new_n344), .A4(new_n262), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n422), .A3(new_n417), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT74), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(new_n417), .A3(new_n422), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n426), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n346), .A2(new_n381), .A3(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n382), .A2(new_n383), .A3(new_n291), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n301), .B1(new_n444), .B2(new_n298), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n281), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT9), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(KEYINPUT72), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT72), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n302), .B2(KEYINPUT9), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n269), .A2(G190), .A3(new_n262), .A4(new_n252), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT73), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n263), .A2(KEYINPUT73), .A3(G190), .A4(new_n269), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n445), .A2(KEYINPUT9), .A3(new_n281), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n270), .A2(G200), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT10), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n451), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n451), .B2(new_n459), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n443), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G244), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n466));
  OAI211_X1 g0266(.A(G238), .B(new_n265), .C1(new_n308), .C2(new_n309), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n466), .B(new_n467), .C1(new_n405), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n246), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n206), .A2(new_n253), .A3(G45), .ZN(new_n471));
  INV_X1    g0271(.A(G250), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n305), .B2(G1), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n327), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT19), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n207), .B1(new_n347), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n406), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n207), .B(G68), .C1(new_n308), .C2(new_n309), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n478), .B1(new_n291), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n301), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n322), .A2(new_n363), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n206), .A2(G33), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n278), .A2(G87), .A3(new_n275), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n474), .B1(new_n469), .B2(new_n246), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n477), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n476), .A2(new_n271), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n486), .A2(new_n301), .B1(new_n363), .B2(new_n322), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n278), .A2(new_n275), .A3(new_n489), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n322), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(new_n339), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OR3_X1    g0301(.A1(new_n275), .A2(KEYINPUT75), .A3(G97), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT75), .B1(new_n275), .B2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n484), .B2(new_n498), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n387), .B2(new_n389), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  AND2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n480), .ZN(new_n509));
  INV_X1    g0309(.A(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(G20), .B1(G77), .B2(new_n295), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n505), .B1(new_n514), .B2(new_n301), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(new_n265), .C1(new_n308), .C2(new_n309), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n246), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT5), .B1(new_n258), .B2(new_n260), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT5), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n206), .B(G45), .C1(new_n525), .C2(G41), .ZN(new_n526));
  OAI211_X1 g0326(.A(G257), .B(new_n327), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n256), .C1(KEYINPUT5), .C2(new_n304), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n523), .A2(G190), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n515), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n529), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n246), .B2(new_n522), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n370), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n495), .B(new_n501), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n524), .A2(new_n526), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n246), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G264), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n472), .A2(G1698), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n308), .B2(new_n309), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT80), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n264), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n543), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n246), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n548), .ZN(new_n552));
  INV_X1    g0352(.A(new_n543), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(new_n553), .A3(new_n550), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n529), .B(new_n540), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  INV_X1    g0356(.A(new_n498), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n275), .A2(new_n558), .A3(G107), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n275), .B2(G107), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n557), .A2(G107), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n510), .A3(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT79), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(new_n567), .A3(new_n568), .A4(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n207), .B(G87), .C1(new_n308), .C2(new_n309), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n264), .A2(new_n576), .A3(new_n207), .A4(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n564), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n578), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n563), .B1(new_n582), .B2(new_n301), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n552), .A2(new_n553), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n549), .A2(new_n550), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n246), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(G190), .A3(new_n529), .A4(new_n540), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n556), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n523), .A2(new_n530), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n295), .A2(G77), .ZN(new_n591));
  INV_X1    g0391(.A(new_n511), .ZN(new_n592));
  XNOR2_X1  g0392(.A(G97), .B(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n507), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n594), .B2(new_n207), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n510), .B1(new_n418), .B2(new_n419), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n301), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n505), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n590), .A2(new_n271), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT76), .B1(new_n534), .B2(new_n339), .ZN(new_n600));
  AND4_X1   g0400(.A1(KEYINPUT76), .A2(new_n523), .A3(new_n339), .A4(new_n530), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n537), .A2(new_n589), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G264), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n604));
  OAI211_X1 g0404(.A(G257), .B(new_n265), .C1(new_n308), .C2(new_n309), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n312), .A2(G303), .A3(new_n313), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n246), .ZN(new_n608));
  OAI211_X1 g0408(.A(G270), .B(new_n327), .C1(new_n524), .C2(new_n526), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n529), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n363), .A2(new_n468), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n278), .A2(G116), .A3(new_n275), .A4(new_n489), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n277), .A2(new_n215), .B1(G20), .B2(new_n468), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n520), .B(new_n207), .C1(G33), .C2(new_n484), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n613), .A2(KEYINPUT20), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT20), .B1(new_n613), .B2(new_n614), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n611), .B(new_n612), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n610), .A2(KEYINPUT21), .A3(G169), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n609), .A2(new_n529), .ZN(new_n619));
  INV_X1    g0419(.A(G179), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n607), .B2(new_n246), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n610), .A2(G169), .A3(new_n617), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT77), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(KEYINPUT77), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n555), .A2(new_n271), .ZN(new_n631));
  INV_X1    g0431(.A(new_n581), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n301), .B1(new_n632), .B2(new_n579), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n562), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n587), .A2(new_n620), .A3(new_n529), .A4(new_n540), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n617), .B1(new_n610), .B2(G200), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT78), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n619), .A2(G190), .A3(new_n608), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(KEYINPUT78), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n630), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n465), .A2(new_n603), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n303), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT84), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n461), .B2(new_n462), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n451), .A2(new_n459), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n451), .A2(new_n459), .A3(new_n460), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(KEYINPUT84), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n379), .A2(new_n380), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n341), .A2(KEYINPUT83), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT83), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n325), .A2(new_n338), .A3(new_n340), .A4(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n653), .B(new_n655), .C1(new_n371), .C2(new_n369), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n441), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(new_n426), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n644), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n501), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n495), .A2(new_n501), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n602), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(G169), .B1(new_n470), .B2(new_n475), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n273), .B(new_n474), .C1(new_n469), .C2(new_n246), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n344), .B(new_n474), .C1(new_n469), .C2(new_n246), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n491), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n499), .A2(new_n666), .B1(new_n668), .B2(new_n477), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT76), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n590), .B2(new_n273), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n534), .A2(KEYINPUT76), .A3(new_n339), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n673), .A4(new_n599), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n660), .B1(new_n663), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n603), .A2(KEYINPUT82), .B1(new_n636), .B2(new_n630), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT82), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n537), .A2(new_n589), .A3(new_n678), .A4(new_n602), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n676), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n659), .B1(new_n465), .B2(new_n680), .ZN(G369));
  AND2_X1   g0481(.A1(new_n630), .A2(new_n641), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT87), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(KEYINPUT85), .B(G343), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT86), .Z(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n617), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n630), .A2(new_n641), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT87), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n630), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n636), .A2(new_n691), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n691), .A2(new_n634), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n589), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n636), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n630), .A2(new_n691), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n210), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n261), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n481), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n213), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n534), .A2(new_n493), .A3(new_n619), .A4(new_n621), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n540), .B1(new_n551), .B2(new_n554), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n619), .A2(new_n493), .A3(new_n621), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n590), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n587), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n610), .A2(new_n339), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n534), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n493), .B(KEYINPUT88), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n555), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n720), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n728), .B2(new_n691), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n556), .A2(new_n583), .A3(new_n588), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n515), .B(new_n531), .C1(new_n370), .C2(new_n534), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n602), .A2(new_n669), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n682), .A3(new_n636), .A4(new_n690), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n716), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n630), .A2(new_n636), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n278), .B1(new_n506), .B2(new_n513), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n534), .A2(G169), .B1(new_n739), .B2(new_n505), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n671), .B2(new_n672), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n536), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n589), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n675), .ZN(new_n744));
  AND4_X1   g0544(.A1(KEYINPUT89), .A2(new_n744), .A3(KEYINPUT29), .A4(new_n690), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n691), .B1(new_n743), .B2(new_n675), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT89), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n680), .B2(new_n691), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n737), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n715), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n709), .A2(new_n350), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G355), .B1(new_n468), .B2(new_n709), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n244), .A2(new_n305), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n709), .A2(new_n264), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G45), .B2(new_n213), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n215), .B1(G20), .B2(new_n271), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n207), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n206), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n710), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n762), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n698), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G50), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n273), .A2(G20), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n344), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n773), .A2(new_n776), .B1(new_n778), .B2(new_n201), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n207), .A2(new_n344), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n273), .A2(new_n370), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(G58), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n484), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n207), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n784), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n370), .A2(G179), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n780), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n406), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n790), .A2(new_n795), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n264), .B1(new_n798), .B2(new_n510), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n273), .A2(new_n370), .A3(new_n790), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n797), .B(new_n799), .C1(new_n801), .C2(G77), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n783), .A2(new_n789), .A3(new_n794), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n776), .A2(new_n804), .B1(new_n805), .B2(new_n787), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT90), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT90), .ZN(new_n808));
  INV_X1    g0608(.A(new_n796), .ZN(new_n809));
  INV_X1    g0609(.A(new_n791), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G303), .A2(new_n809), .B1(new_n810), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n350), .C1(new_n812), .C2(new_n798), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G322), .B2(new_n782), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n777), .A2(new_n815), .B1(new_n801), .B2(G311), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n807), .A2(new_n808), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n770), .B(new_n772), .C1(new_n763), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n700), .A2(new_n769), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n698), .A2(G330), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  OAI21_X1  g0624(.A(KEYINPUT82), .B1(new_n732), .B2(new_n734), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(new_n679), .A3(new_n738), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n691), .B1(new_n826), .B2(new_n675), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n690), .A2(new_n324), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n653), .A2(new_n655), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n345), .B(new_n341), .C1(new_n324), .C2(new_n690), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n827), .B(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n737), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n769), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(new_n769), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n763), .A2(new_n760), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT91), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n836), .B1(new_n839), .B2(new_n202), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G283), .A2(new_n777), .B1(new_n775), .B2(G303), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n468), .B2(new_n800), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT92), .ZN(new_n843));
  INV_X1    g0643(.A(new_n798), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G87), .A2(new_n844), .B1(new_n810), .B2(G311), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(new_n350), .C1(new_n510), .C2(new_n796), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n788), .B(new_n846), .C1(G294), .C2(new_n782), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT93), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G143), .A2(new_n782), .B1(new_n801), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n776), .B2(new_n851), .C1(new_n294), .C2(new_n778), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n264), .B1(new_n796), .B2(new_n773), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n798), .A2(new_n201), .B1(new_n791), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(G58), .C2(new_n786), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n848), .A2(KEYINPUT93), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n849), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n763), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n840), .B1(new_n761), .B2(new_n831), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n835), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  OR2_X1    g0666(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(G116), .A3(new_n216), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI211_X1 g0670(.A(new_n214), .B(G77), .C1(new_n285), .C2(new_n201), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n773), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n206), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n731), .A2(new_n736), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n691), .A2(new_n380), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n381), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n380), .B(new_n691), .C1(new_n379), .C2(new_n372), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n831), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n416), .A2(new_n423), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n423), .A2(new_n687), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n435), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .A4(new_n435), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n882), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n426), .B2(new_n441), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n880), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n737), .A2(new_n464), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT96), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n464), .A2(new_n875), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n879), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n827), .A2(new_n831), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n691), .A2(new_n341), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n887), .A2(new_n889), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT94), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n890), .B2(new_n891), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n913), .A2(KEYINPUT94), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT95), .Z(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n914), .A3(new_n917), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n379), .A2(new_n380), .A3(new_n690), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n687), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n426), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n912), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n751), .B(new_n464), .C1(new_n747), .C2(new_n745), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n659), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n926), .B(new_n928), .Z(new_n929));
  OAI22_X1  g0729(.A1(new_n901), .A2(new_n929), .B1(new_n206), .B2(new_n766), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n901), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n874), .B1(new_n930), .B2(new_n931), .ZN(G367));
  INV_X1    g0732(.A(new_n757), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n764), .B1(new_n210), .B2(new_n322), .C1(new_n933), .C2(new_n234), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n510), .B2(new_n787), .ZN(new_n936));
  INV_X1    g0736(.A(G317), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n350), .B1(new_n791), .B2(new_n937), .C1(new_n484), .C2(new_n798), .ZN(new_n938));
  INV_X1    g0738(.A(G303), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n781), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT46), .B1(new_n809), .B2(G116), .ZN(new_n941));
  NOR4_X1   g0741(.A1(new_n936), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n777), .A2(G294), .B1(new_n801), .B2(G283), .ZN(new_n943));
  INV_X1    g0743(.A(G311), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n776), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G58), .A2(new_n809), .B1(new_n844), .B2(G77), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n350), .B1(new_n810), .B2(G137), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n201), .C2(new_n787), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G50), .A2(new_n801), .B1(new_n782), .B2(G150), .ZN(new_n949));
  INV_X1    g0749(.A(G143), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n949), .B1(new_n776), .B2(new_n950), .C1(new_n792), .C2(new_n778), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n945), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT47), .Z(new_n953));
  OAI211_X1 g0753(.A(new_n769), .B(new_n934), .C1(new_n953), .C2(new_n863), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n691), .A2(new_n491), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n662), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n771), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n704), .A2(new_n706), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT103), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n699), .B(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n704), .A2(new_n706), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n752), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n707), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n741), .A2(new_n690), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n733), .B1(new_n690), .B2(new_n515), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n975), .A2(new_n602), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n971), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n707), .A2(new_n977), .A3(new_n970), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n707), .A2(new_n977), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(KEYINPUT102), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n705), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n987), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT102), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n969), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n986), .A2(new_n705), .A3(new_n987), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT104), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n986), .A2(KEYINPUT104), .A3(new_n705), .A4(new_n987), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n961), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n989), .A3(new_n988), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n969), .ZN(new_n1002));
  AND4_X1   g0802(.A1(new_n961), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n752), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n710), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n768), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n704), .A2(new_n706), .A3(new_n977), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT97), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT42), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n631), .A2(new_n634), .A3(new_n635), .A4(new_n733), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n691), .B1(new_n1013), .B2(new_n602), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT98), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(KEYINPUT98), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n705), .A2(new_n978), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT43), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1016), .A2(new_n1017), .A3(new_n1021), .A4(new_n956), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1020), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n960), .B1(new_n1008), .B2(new_n1026), .ZN(G387));
  XNOR2_X1  g0827(.A(new_n965), .B(new_n966), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n704), .A2(new_n771), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n754), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(new_n712), .B1(G107), .B2(new_n210), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT106), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n283), .A2(G50), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT50), .Z(new_n1034));
  NAND3_X1  g0834(.A1(new_n712), .A2(new_n305), .A3(new_n240), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n757), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT107), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n231), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(G45), .B1(KEYINPUT107), .B2(new_n1036), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1032), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n764), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n769), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n776), .A2(new_n792), .B1(new_n201), .B2(new_n800), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G50), .B2(new_n782), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n382), .A2(new_n383), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n777), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n787), .A2(new_n322), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n264), .B1(new_n798), .B2(new_n484), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n796), .A2(new_n202), .B1(new_n791), .B2(new_n294), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1044), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n264), .B1(new_n810), .B2(G326), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n787), .A2(new_n812), .B1(new_n796), .B2(new_n805), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G303), .A2(new_n801), .B1(new_n782), .B2(G317), .ZN(new_n1054));
  INV_X1    g0854(.A(G322), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1054), .B1(new_n776), .B2(new_n1055), .C1(new_n944), .C2(new_n778), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT49), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT108), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1052), .B1(new_n468), .B2(new_n798), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1060), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT108), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1051), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1042), .B1(new_n1065), .B2(new_n763), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1028), .A2(new_n768), .B1(new_n1029), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n969), .A2(new_n710), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1028), .A2(new_n752), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  OAI21_X1  g0870(.A(new_n764), .B1(new_n484), .B2(new_n210), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n757), .B2(new_n238), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n836), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n264), .B1(new_n798), .B2(new_n406), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n787), .A2(new_n202), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT109), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n796), .A2(new_n201), .B1(new_n791), .B2(new_n950), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1074), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1077), .A2(new_n1076), .B1(new_n800), .B2(new_n283), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G50), .B2(new_n777), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n775), .A2(G150), .B1(new_n782), .B2(G159), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1078), .B(new_n1080), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n775), .A2(G317), .B1(new_n782), .B2(G311), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT110), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G283), .A2(new_n809), .B1(new_n810), .B2(G322), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n264), .B1(new_n844), .B2(G107), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n468), .C2(new_n787), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n778), .A2(new_n939), .B1(new_n805), .B2(new_n800), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1086), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1073), .B1(new_n1096), .B2(new_n863), .C1(new_n771), .C2(new_n977), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n991), .A2(new_n989), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n999), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n767), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n994), .A2(new_n961), .A3(new_n999), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n988), .A2(new_n989), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT102), .B1(new_n986), .B2(new_n987), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n752), .B(new_n1028), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n997), .A2(new_n998), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT105), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n711), .B1(new_n1099), .B2(new_n969), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1100), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  OR3_X1    g0910(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n294), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT53), .B1(new_n796), .B2(new_n294), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n792), .C2(new_n787), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n350), .B1(new_n810), .B2(G125), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n773), .B2(new_n798), .C1(new_n778), .C2(new_n851), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT115), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1113), .B(new_n1115), .C1(new_n801), .C2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n775), .A2(G128), .B1(new_n782), .B2(G132), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT116), .Z(new_n1120));
  OAI22_X1  g0920(.A1(new_n776), .A2(new_n812), .B1(new_n468), .B2(new_n781), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n798), .A2(new_n201), .B1(new_n791), .B2(new_n805), .ZN(new_n1122));
  OR4_X1    g0922(.A1(new_n264), .A2(new_n1075), .A3(new_n797), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n778), .A2(new_n510), .B1(new_n484), .B2(new_n800), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1121), .B(new_n1123), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1125), .A2(new_n1124), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1118), .A2(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n769), .B1(new_n1045), .B2(new_n838), .C1(new_n1128), .C2(new_n863), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n919), .A2(new_n920), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n760), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n728), .A2(new_n691), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT31), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n603), .A2(new_n642), .A3(new_n691), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n831), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n902), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n892), .A2(new_n922), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(KEYINPUT111), .B(new_n904), .C1(new_n746), .C2(new_n831), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT111), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n744), .A2(new_n690), .A3(new_n831), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n905), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1141), .B1(new_n1146), .B2(new_n879), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n829), .A2(new_n830), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n691), .B(new_n1148), .C1(new_n826), .C2(new_n675), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n879), .B1(new_n1149), .B2(new_n904), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1150), .A2(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1139), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1130), .B1(new_n906), .B2(new_n922), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1144), .A2(new_n905), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT111), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1144), .A2(new_n1143), .A3(new_n905), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n879), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1140), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n737), .A2(new_n831), .A3(new_n879), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1153), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1131), .B1(new_n1162), .B2(new_n768), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n464), .B1(new_n827), .B2(KEYINPUT29), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n659), .B(new_n897), .C1(new_n748), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT112), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT112), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n927), .A2(new_n1167), .A3(new_n659), .A4(new_n897), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n903), .A2(new_n905), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n879), .B1(new_n737), .B2(new_n831), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1169), .B1(new_n1139), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1138), .A2(new_n902), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1159), .B(new_n1172), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT113), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1166), .A2(new_n1168), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1166), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT113), .ZN(new_n1178));
  AOI211_X1 g0978(.A(KEYINPUT114), .B(new_n1161), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT114), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1176), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1162), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n710), .B1(new_n1181), .B2(new_n1162), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1163), .B1(new_n1183), .B2(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(new_n1162), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT114), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1181), .A2(new_n1180), .A3(new_n1162), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n651), .A2(new_n303), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n446), .A3(new_n687), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n651), .B(new_n303), .C1(new_n302), .C2(new_n924), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n896), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n926), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n896), .A2(new_n1198), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n926), .B1(new_n1204), .B2(new_n1199), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1186), .B1(new_n1191), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1187), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1186), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n711), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1198), .A2(new_n760), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n777), .A2(G97), .B1(new_n782), .B2(G107), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n468), .B2(new_n776), .C1(new_n322), .C2(new_n800), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n787), .A2(new_n201), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n796), .A2(new_n202), .B1(new_n791), .B2(new_n812), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n350), .B(new_n304), .C1(new_n798), .C2(new_n285), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT118), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n787), .A2(new_n294), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n775), .B2(G125), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n777), .A2(G132), .B1(new_n801), .B2(G137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1117), .A2(new_n809), .B1(new_n782), .B2(G128), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT119), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1225), .B(new_n1226), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n405), .B(new_n257), .C1(new_n798), .C2(new_n792), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G124), .B2(new_n810), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n773), .B1(G33), .B2(G41), .C1(new_n261), .C2(new_n264), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1223), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n763), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n836), .B1(new_n839), .B2(new_n773), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1214), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1206), .B2(new_n768), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1213), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT120), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n902), .A2(new_n760), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n769), .B1(new_n838), .B2(G68), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1047), .B1(G283), .B2(new_n782), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT121), .Z(new_n1250));
  OAI21_X1  g1050(.A(new_n350), .B1(new_n798), .B2(new_n202), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n796), .A2(new_n484), .B1(new_n791), .B2(new_n939), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n777), .C2(G116), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n775), .A2(G294), .B1(new_n801), .B2(G107), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n775), .A2(G132), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT122), .Z(new_n1257));
  OAI21_X1  g1057(.A(new_n264), .B1(new_n798), .B2(new_n285), .ZN(new_n1258));
  INV_X1    g1058(.A(G128), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n796), .A2(new_n792), .B1(new_n791), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G50), .C2(new_n786), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n777), .A2(new_n1117), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G137), .A2(new_n782), .B1(new_n801), .B2(G150), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1255), .B1(new_n1257), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1248), .B1(new_n1265), .B2(new_n763), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1174), .A2(new_n768), .B1(new_n1247), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1181), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1209), .A2(new_n1174), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1271), .B2(new_n1006), .ZN(G381));
  INV_X1    g1072(.A(G375), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n752), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n767), .B1(new_n1275), .B2(new_n1006), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n959), .B1(new_n1276), .B2(new_n1025), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1278));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1109), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n1277), .A3(new_n1280), .ZN(G407));
  INV_X1    g1081(.A(G213), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n688), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(new_n1279), .A3(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(G407), .A2(new_n1284), .A3(G213), .ZN(G409));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1206), .A2(KEYINPUT124), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n767), .B1(new_n1206), .B2(KEYINPUT124), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1243), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1210), .A2(new_n1007), .A3(new_n1206), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G378), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1201), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1204), .A2(new_n1199), .A3(new_n926), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT57), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n710), .B1(new_n1191), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1206), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G378), .B(new_n1244), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT123), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1213), .A2(new_n1299), .A3(G378), .A4(new_n1244), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1291), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1271), .A2(KEYINPUT60), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1302), .B(new_n710), .C1(KEYINPUT60), .C2(new_n1269), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1267), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n865), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(G384), .A3(new_n1267), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1301), .A2(new_n1283), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1286), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1291), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1244), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1299), .B1(new_n1314), .B2(G378), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1311), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1283), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1283), .A2(G2897), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1307), .B(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1307), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1317), .A3(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1310), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(G393), .B(new_n823), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1276), .A2(new_n1025), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G390), .B1(new_n1328), .B2(new_n960), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n959), .B(new_n1109), .C1(new_n1276), .C2(new_n1025), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1327), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(new_n1109), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1277), .A2(G390), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1326), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1325), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1335), .B1(new_n1323), .B2(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1338), .B(new_n1321), .C1(new_n1337), .C2(new_n1323), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(G405));
  NAND3_X1  g1140(.A1(new_n1335), .A2(KEYINPUT126), .A3(new_n1322), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1322), .A2(KEYINPUT126), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1331), .A2(new_n1334), .A3(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(G375), .A2(new_n1279), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT127), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1345), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1344), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT127), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1345), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1353));
  AOI22_X1  g1153(.A1(new_n1352), .A2(new_n1353), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1350), .A2(new_n1354), .ZN(G402));
endmodule


