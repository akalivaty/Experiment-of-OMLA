//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT0), .A4(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n201), .B2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(KEYINPUT66), .A3(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n202), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n210), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n198), .A2(new_n208), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n222), .A3(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n189), .A2(G137), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n191), .A2(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n197), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(KEYINPUT2), .A2(G113), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(KEYINPUT2), .B2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT68), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n233), .C1(new_n235), .C2(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n200), .A2(new_n202), .A3(G128), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n222), .A2(new_n244), .B1(new_n214), .B2(new_n220), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n197), .A2(new_n227), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n224), .A2(new_n228), .A3(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n218), .A3(new_n249), .A4(KEYINPUT30), .ZN(new_n250));
  AND4_X1   g064(.A1(KEYINPUT70), .A2(new_n232), .A3(new_n243), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n243), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n230), .B2(new_n231), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT70), .B1(new_n253), .B2(new_n250), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT31), .ZN(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  INV_X1    g072(.A(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n260), .B(new_n261), .Z(new_n262));
  NAND4_X1  g076(.A1(new_n247), .A2(new_n252), .A3(new_n218), .A4(new_n249), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n255), .A2(new_n256), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n232), .A2(new_n243), .A3(new_n250), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n250), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n262), .A3(new_n263), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n230), .A2(new_n243), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n230), .B2(new_n243), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n262), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n273), .A2(new_n263), .ZN(new_n283));
  INV_X1    g097(.A(new_n272), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n278), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n262), .ZN(new_n289));
  INV_X1    g103(.A(new_n262), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n255), .A2(new_n290), .A3(new_n263), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n247), .A2(new_n218), .A3(new_n249), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n243), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT73), .A3(new_n263), .ZN(new_n297));
  OR3_X1    g111(.A1(new_n295), .A2(KEYINPUT73), .A3(new_n243), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT28), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n278), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G472), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n288), .A2(new_n290), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n264), .A3(new_n270), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G128), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n308), .A2(KEYINPUT23), .A3(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(G119), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT23), .B1(new_n308), .B2(G119), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G110), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G110), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G128), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(KEYINPUT75), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n308), .B2(G119), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n310), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT24), .B(G110), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(KEYINPUT78), .A2(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(KEYINPUT78), .A2(G125), .ZN(new_n329));
  OAI21_X1  g143(.A(G140), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n331), .A3(G125), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(KEYINPUT16), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n328), .A2(new_n329), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT16), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n331), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n339), .A3(G146), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(G146), .B1(new_n336), .B2(new_n339), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n320), .B(new_n327), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n325), .A2(new_n326), .B1(new_n317), .B2(G110), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n331), .A2(G125), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n199), .A3(new_n332), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n343), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n343), .B2(new_n347), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n356), .A2(new_n294), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n294), .A3(new_n353), .A4(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n358), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n294), .B2(G234), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n307), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(G104), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n377), .A2(G107), .B1(KEYINPUT82), .B2(KEYINPUT3), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n377), .A2(G107), .B1(KEYINPUT82), .B2(KEYINPUT3), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .A4(new_n259), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n375), .A2(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n377), .A2(G107), .ZN(new_n382));
  OAI21_X1  g196(.A(G101), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n221), .B2(new_n223), .ZN(new_n386));
  AND4_X1   g200(.A1(new_n222), .A2(new_n200), .A3(new_n202), .A4(G128), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n219), .A2(G128), .B1(new_n200), .B2(new_n202), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n380), .B(new_n383), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n384), .A2(new_n386), .B1(new_n389), .B2(new_n385), .ZN(new_n390));
  INV_X1    g204(.A(new_n198), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n396), .A3(new_n208), .A4(new_n217), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n389), .B1(new_n384), .B2(new_n224), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n399), .A2(KEYINPUT12), .A3(new_n198), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT12), .B1(new_n399), .B2(new_n198), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  INV_X1    g219(.A(G227), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G953), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n405), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n398), .B(KEYINPUT83), .C1(new_n400), .C2(new_n401), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n409), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n391), .B1(new_n390), .B2(new_n397), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT84), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n408), .B1(new_n402), .B2(new_n403), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n421), .A2(new_n410), .B1(new_n415), .B2(new_n413), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(G469), .C1(new_n422), .C2(G902), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n409), .B1(new_n412), .B2(new_n414), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n398), .B(new_n408), .C1(new_n400), .C2(new_n401), .ZN(new_n425));
  AOI211_X1 g239(.A(G469), .B(new_n293), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT9), .B(G234), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT81), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n394), .A2(new_n243), .A3(new_n396), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n321), .A2(G116), .ZN(new_n441));
  INV_X1    g255(.A(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G119), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT5), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(G113), .C1(KEYINPUT5), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n242), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n380), .A2(new_n383), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n384), .A2(KEYINPUT85), .A3(new_n242), .A4(new_n445), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n439), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n456), .A3(new_n452), .ZN(new_n457));
  INV_X1    g271(.A(new_n337), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n208), .B2(new_n217), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n224), .A2(new_n337), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n461), .B(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n455), .A2(new_n457), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G902), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n459), .A2(new_n460), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n471));
  OAI221_X1 g285(.A(new_n471), .B1(new_n468), .B2(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n472));
  INV_X1    g286(.A(new_n459), .ZN(new_n473));
  INV_X1    g287(.A(new_n460), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n468), .B1(new_n463), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(KEYINPUT87), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n474), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n451), .B(KEYINPUT8), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n446), .A2(new_n447), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n446), .A2(new_n447), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n470), .A2(new_n472), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n454), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n467), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n438), .B1(new_n466), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n455), .A2(new_n457), .A3(new_n465), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n478), .A2(new_n482), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(new_n454), .A3(new_n470), .A4(new_n472), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n487), .A2(new_n489), .A3(new_n467), .A4(new_n437), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n436), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n349), .A2(G952), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(G234), .B2(G237), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n349), .B(new_n294), .C1(G234), .C2(G237), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT21), .B(G898), .Z(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(G143), .B1(new_n257), .B2(G214), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n257), .A2(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n201), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n196), .A3(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  MUX2_X1   g321(.A(new_n507), .B(new_n503), .S(KEYINPUT17), .Z(new_n508));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n341), .B2(new_n342), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n336), .A2(new_n339), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n199), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT90), .A3(new_n340), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n505), .A2(new_n500), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G146), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n346), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G113), .B(G122), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT88), .B(G104), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n514), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n514), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n467), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G475), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n507), .A2(new_n340), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n345), .A2(new_n332), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT19), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n518), .B2(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n199), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n532), .A2(new_n536), .B1(new_n520), .B2(new_n517), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n530), .B1(new_n537), .B2(new_n524), .ZN(new_n538));
  AOI211_X1 g352(.A(G146), .B(new_n534), .C1(new_n518), .C2(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n521), .B1(new_n539), .B2(new_n531), .ZN(new_n540));
  INV_X1    g354(.A(new_n524), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT89), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n525), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n529), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n442), .A2(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT91), .B(G122), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n442), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n375), .ZN(new_n553));
  OAI211_X1 g367(.A(G107), .B(new_n550), .C1(new_n551), .C2(new_n442), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT14), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G122), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n556), .B1(new_n561), .B2(G116), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  XNOR2_X1  g377(.A(G128), .B(G143), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G134), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n308), .A2(G143), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n201), .A2(G128), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n189), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n555), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n308), .A2(G143), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT92), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT13), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(G134), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n568), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n564), .A2(G134), .A3(new_n573), .A4(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n562), .A2(G107), .A3(new_n568), .A4(new_n565), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n553), .A4(new_n554), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n429), .A2(G217), .A3(new_n349), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n570), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n570), .B2(new_n581), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n549), .B(new_n294), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT15), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(G478), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n570), .A2(new_n581), .ZN(new_n588));
  INV_X1    g402(.A(new_n582), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n570), .A2(new_n581), .A3(new_n582), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n586), .A2(G478), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n549), .A3(new_n294), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n499), .A2(new_n548), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT80), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n307), .A2(new_n598), .A3(new_n371), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n373), .A2(new_n434), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n305), .A2(new_n294), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(new_n428), .A3(new_n433), .A4(new_n280), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n583), .B2(new_n584), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n590), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n294), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G478), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n611), .A3(new_n294), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n609), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n548), .ZN(new_n616));
  NOR4_X1   g430(.A1(new_n604), .A2(new_n499), .A3(new_n370), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n305), .B2(new_n294), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n187), .B2(new_n305), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n595), .B(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n499), .A2(new_n548), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n434), .A2(new_n624), .A3(new_n627), .A4(new_n371), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n343), .A2(new_n347), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n343), .B2(new_n347), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT98), .B1(new_n634), .B2(new_n368), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  INV_X1    g450(.A(new_n368), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n632), .A2(new_n633), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n367), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n434), .A2(new_n624), .A3(new_n597), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n640), .B(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT32), .B1(new_n305), .B2(new_n187), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n649), .B2(new_n303), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n428), .A2(new_n433), .A3(new_n491), .ZN(new_n651));
  INV_X1    g465(.A(new_n547), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n652), .A2(new_n653), .B1(G475), .B2(new_n528), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n493), .B1(new_n495), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n596), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n656), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n434), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n548), .B(new_n596), .C1(new_n663), .C2(KEYINPUT40), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(KEYINPUT40), .B2(new_n663), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n367), .A2(new_n639), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n290), .B1(new_n255), .B2(new_n263), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n297), .A2(new_n298), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n467), .B1(new_n668), .B2(new_n262), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n282), .A2(new_n306), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n486), .A2(new_n490), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT38), .Z(new_n674));
  NOR3_X1   g488(.A1(new_n672), .A2(new_n436), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n665), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  INV_X1    g491(.A(new_n651), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n609), .A2(new_n612), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT95), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n548), .A2(new_n680), .A3(new_n681), .A4(new_n657), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n678), .A2(new_n307), .A3(new_n641), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  NOR2_X1   g499(.A1(new_n616), .A2(new_n499), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n424), .A2(new_n425), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n418), .B1(new_n687), .B2(new_n294), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n426), .A3(new_n432), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n307), .A3(new_n371), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n307), .A2(new_n627), .A3(new_n371), .A4(new_n689), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND4_X1  g509(.A1(new_n307), .A2(new_n597), .A3(new_n641), .A4(new_n689), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND3_X1  g511(.A1(new_n299), .A2(KEYINPUT101), .A3(new_n278), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n290), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT101), .B1(new_n299), .B2(new_n278), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n264), .B(new_n270), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n623), .B1(new_n187), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n499), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n596), .A2(new_n548), .A3(new_n689), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n371), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  AND2_X1   g520(.A1(new_n491), .A2(new_n689), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n187), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n603), .A2(new_n707), .A3(new_n640), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n682), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n615), .A2(KEYINPUT102), .A3(new_n548), .A4(new_n657), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n427), .B1(new_n417), .B2(new_n418), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n673), .A2(new_n432), .A3(new_n436), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n307), .A2(new_n371), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n370), .B1(new_n649), .B2(new_n303), .ZN(new_n722));
  INV_X1    g536(.A(new_n717), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n711), .B2(new_n712), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT42), .A4(new_n719), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  OR3_X1    g541(.A1(new_n720), .A2(new_n658), .A3(new_n723), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  OR2_X1    g543(.A1(new_n422), .A2(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n422), .A2(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(G469), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(G469), .A2(G902), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n427), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT103), .B1(new_n735), .B2(new_n427), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n433), .A3(new_n662), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n615), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n548), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(KEYINPUT43), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n624), .A2(new_n666), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT44), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n673), .A2(new_n436), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n751), .A2(new_n753), .A3(KEYINPUT44), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n740), .A2(KEYINPUT104), .A3(new_n433), .A4(new_n662), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n743), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  NAND3_X1  g575(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n433), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n739), .B2(new_n432), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n307), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n370), .A3(new_n683), .A4(new_n755), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  NAND4_X1  g581(.A1(new_n690), .A2(new_n694), .A3(new_n696), .A4(new_n705), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n595), .B(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n499), .A2(new_n548), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n434), .A2(new_n624), .A3(new_n771), .A4(new_n371), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n642), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n642), .A2(new_n772), .A3(KEYINPUT110), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n768), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n307), .A2(new_n598), .A3(new_n371), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n598), .B1(new_n307), .B2(new_n371), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n434), .A2(new_n597), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(KEYINPUT108), .A3(new_n617), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  INV_X1    g597(.A(new_n617), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n600), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n777), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n702), .A2(new_n640), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n724), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n307), .A2(new_n428), .A3(new_n641), .A4(new_n657), .ZN(new_n790));
  INV_X1    g604(.A(new_n770), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n548), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n719), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n726), .A3(new_n728), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n433), .A2(new_n666), .A3(new_n657), .A4(new_n717), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n596), .A2(new_n491), .A3(new_n548), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n671), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n671), .A2(new_n797), .A3(KEYINPUT111), .A4(new_n798), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n660), .A2(new_n684), .A3(new_n714), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n796), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n802), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n651), .A2(new_n682), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n650), .A2(new_n807), .B1(new_n709), .B2(new_n713), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n808), .A3(KEYINPUT52), .A4(new_n660), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n805), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n814), .B(new_n796), .C1(new_n803), .C2(new_n804), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n795), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n812), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(new_n719), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n688), .A2(new_n426), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n494), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(new_n672), .A3(new_n371), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n548), .A3(new_n615), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n795), .A2(new_n818), .A3(KEYINPUT53), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n726), .A2(new_n728), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n307), .A2(new_n428), .A3(new_n641), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n654), .A3(new_n657), .A4(new_n770), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n824), .B1(new_n835), .B2(new_n788), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT108), .B1(new_n781), .B2(new_n617), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n600), .A2(new_n784), .A3(new_n783), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n810), .A2(new_n837), .A3(new_n777), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n820), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n823), .A2(new_n829), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n493), .A2(new_n751), .A3(new_n371), .A4(new_n702), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n689), .A2(new_n436), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT116), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n674), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(KEYINPUT50), .A3(new_n674), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n762), .A2(new_n764), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n826), .A2(new_n433), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n755), .B(new_n847), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n828), .A2(new_n654), .A3(new_n744), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n751), .A2(new_n827), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n787), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n857), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT51), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n492), .B1(new_n862), .B2(new_n864), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n847), .A2(new_n707), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n722), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT48), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n846), .A2(new_n870), .B1(G952), .B2(G953), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n674), .A2(new_n371), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n432), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n435), .A3(new_n672), .A4(new_n745), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(G75));
  AOI21_X1  g691(.A(new_n294), .B1(new_n830), .B2(new_n842), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n438), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n878), .B2(new_n438), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n455), .A2(new_n457), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n465), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT55), .Z(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n881), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n349), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n879), .A2(new_n882), .A3(new_n880), .A4(new_n886), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT119), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n888), .A2(new_n894), .A3(new_n890), .A4(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n733), .A2(KEYINPUT57), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n733), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g712(.A(new_n843), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n832), .B1(new_n830), .B2(new_n842), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n897), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n687), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n732), .B(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n878), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n889), .B1(new_n902), .B2(new_n904), .ZN(G54));
  AND3_X1   g719(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(new_n543), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n543), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n889), .ZN(G60));
  NAND2_X1  g723(.A1(new_n606), .A2(new_n607), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT59), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(new_n913), .C1(new_n899), .C2(new_n900), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n916), .B(new_n812), .C1(new_n811), .C2(new_n821), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n845), .A2(new_n844), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n889), .B(new_n915), .C1(new_n919), .C2(new_n910), .ZN(G63));
  NAND2_X1  g734(.A1(new_n830), .A2(new_n842), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n365), .A2(new_n467), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n356), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(KEYINPUT122), .A3(new_n924), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT122), .B1(new_n921), .B2(new_n924), .ZN(new_n931));
  INV_X1    g745(.A(new_n924), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n926), .B(new_n932), .C1(new_n830), .C2(new_n842), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n634), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n930), .A2(new_n934), .A3(new_n890), .A4(new_n936), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G66));
  AOI21_X1  g753(.A(new_n349), .B1(new_n497), .B2(G224), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n786), .B2(new_n349), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT124), .ZN(new_n942));
  INV_X1    g756(.A(G898), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n884), .B1(new_n943), .B2(G953), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G69));
  NAND2_X1  g759(.A1(new_n232), .A2(new_n250), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n535), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n804), .B(KEYINPUT126), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n676), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT62), .Z(new_n952));
  NOR2_X1   g766(.A1(new_n663), .A2(new_n756), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n616), .B1(new_n548), .B2(new_n770), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n953), .A2(new_n373), .A3(new_n599), .A4(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n952), .A2(new_n760), .A3(new_n766), .A4(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n956), .B2(new_n349), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n766), .A2(new_n760), .A3(new_n950), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n743), .A2(new_n722), .A3(new_n759), .A4(new_n798), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n726), .A3(new_n728), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n349), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n655), .A2(G953), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT127), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n948), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n349), .B1(G227), .B2(G900), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n957), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n957), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n956), .B2(new_n786), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n889), .B1(new_n971), .B2(new_n667), .ZN(new_n972));
  INV_X1    g786(.A(new_n291), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n958), .A2(new_n960), .A3(new_n786), .ZN(new_n974));
  INV_X1    g788(.A(new_n970), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n973), .A2(new_n667), .A3(new_n975), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n822), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n972), .A2(new_n976), .A3(new_n978), .ZN(G57));
endmodule


