//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n210), .B(new_n211), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(G113gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G120gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT64), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n230), .A2(new_n234), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n228), .ZN(new_n240));
  OR2_X1    g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n226), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n229), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT66), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n248), .A2(new_n241), .A3(new_n226), .A4(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n239), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n246), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(G190gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(KEYINPUT28), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n255), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n254), .A2(new_n255), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(KEYINPUT28), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n238), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n263));
  OR3_X1    g062(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n225), .B1(new_n253), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n244), .A2(new_n245), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n239), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n245), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n224), .A3(new_n267), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n204), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(new_n204), .A3(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT34), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n278), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(KEYINPUT32), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(new_n277), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G71gat), .B(G99gat), .Z(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT73), .B(G15gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n291));
  INV_X1    g090(.A(G43gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n290), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n278), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT33), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n282), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n282), .B2(new_n287), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT36), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n280), .A2(new_n281), .A3(new_n277), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n287), .A3(new_n297), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT36), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT0), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(G57gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G85gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G141gat), .B(G148gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n318), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT77), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n224), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n324), .A2(new_n334), .B1(G155gat), .B2(G162gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n315), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(new_n325), .B1(new_n213), .B2(new_n223), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n314), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT4), .B1(new_n332), .B2(new_n224), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n317), .A2(new_n318), .B1(new_n321), .B2(new_n323), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n335), .B2(new_n337), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n213), .A4(new_n223), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n224), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n313), .A3(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n341), .A2(new_n352), .A3(KEYINPUT79), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n341), .B1(KEYINPUT79), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n312), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT6), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(KEYINPUT79), .ZN(new_n357));
  INV_X1    g156(.A(new_n341), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n352), .A3(KEYINPUT79), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n311), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n353), .A2(new_n354), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n311), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  INV_X1    g165(.A(G197gat), .ZN(new_n367));
  INV_X1    g166(.A(G204gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT22), .ZN(new_n371));
  NAND2_X1  g170(.A1(G211gat), .A2(G218gat), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n369), .A2(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  NOR2_X1   g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT74), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G211gat), .ZN(new_n377));
  INV_X1    g176(.A(G218gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n372), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n373), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n369), .A2(new_n370), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n371), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n376), .A2(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n366), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(new_n381), .ZN(new_n387));
  INV_X1    g186(.A(new_n373), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n376), .A3(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n275), .A2(new_n267), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n275), .B2(new_n267), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n392), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n253), .B2(new_n268), .ZN(new_n400));
  INV_X1    g199(.A(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n275), .A2(new_n267), .A3(new_n393), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G64gat), .ZN(new_n405));
  INV_X1    g204(.A(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n399), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n399), .B2(new_n403), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT76), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n394), .A2(new_n398), .A3(new_n392), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT30), .A4(new_n408), .ZN(new_n418));
  AND4_X1   g217(.A1(new_n365), .A2(new_n412), .A3(new_n413), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n395), .B1(new_n332), .B2(KEYINPUT3), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n349), .A2(new_n422), .A3(new_n395), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(new_n392), .ZN(new_n424));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n395), .B1(new_n382), .B2(new_n385), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n344), .B1(new_n427), .B2(new_n348), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n392), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT81), .B1(new_n392), .B2(new_n420), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n431), .A2(new_n432), .A3(new_n428), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  INV_X1    g233(.A(G22gat), .ZN(new_n435));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT31), .ZN(new_n437));
  INV_X1    g236(.A(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n434), .A2(new_n435), .B1(KEYINPUT80), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n392), .A2(new_n420), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n392), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n429), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n425), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(G22gat), .A3(new_n430), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n446), .B(new_n430), .C1(KEYINPUT83), .C2(new_n435), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n440), .A2(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n439), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n419), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT84), .B1(new_n307), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n412), .A2(new_n418), .A3(new_n413), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n347), .A2(new_n351), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n314), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n333), .A2(new_n339), .A3(new_n314), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n311), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n314), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n463), .A2(KEYINPUT87), .A3(KEYINPUT40), .A4(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n344), .A2(new_n348), .B1(new_n213), .B2(new_n223), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n342), .A2(new_n346), .B1(new_n467), .B2(new_n350), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT39), .B(new_n462), .C1(new_n468), .C2(new_n313), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(new_n312), .A3(KEYINPUT40), .A4(new_n465), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n312), .A3(new_n465), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT86), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(KEYINPUT86), .A3(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n473), .B(new_n361), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n457), .B1(new_n458), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n399), .A2(new_n481), .A3(new_n403), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n407), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n399), .B2(new_n403), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT38), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n483), .A2(KEYINPUT38), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n403), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(KEYINPUT37), .C1(KEYINPUT89), .C2(new_n399), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n362), .A2(new_n364), .A3(new_n409), .ZN(new_n492));
  OAI211_X1 g291(.A(KEYINPUT90), .B(KEYINPUT38), .C1(new_n483), .C2(new_n484), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n487), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n412), .A2(new_n418), .A3(new_n413), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n475), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n498), .A2(new_n477), .B1(new_n363), .B2(new_n311), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n495), .A2(new_n499), .A3(KEYINPUT88), .A4(new_n473), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n494), .A3(new_n454), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n304), .A2(KEYINPUT36), .A3(new_n305), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n434), .A2(new_n435), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n447), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n450), .A2(new_n451), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n504), .A2(new_n447), .A3(new_n505), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n508), .A2(new_n439), .B1(new_n509), .B2(KEYINPUT80), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n365), .A2(new_n412), .A3(new_n413), .A4(new_n418), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n502), .A2(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n456), .A2(new_n501), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n419), .A2(new_n454), .A3(new_n305), .A4(new_n304), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(KEYINPUT92), .A3(new_n523), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n528), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n438), .A2(G43gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n292), .A2(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n535), .A2(KEYINPUT96), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(KEYINPUT96), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n538), .B(new_n539), .C1(G43gat), .C2(new_n438), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n540), .B2(new_n536), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n545), .A2(KEYINPUT94), .A3(new_n546), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n546), .B2(KEYINPUT94), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n537), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n533), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n554), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT17), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n557), .B2(new_n533), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT97), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n533), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n556), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n559), .B(KEYINPUT13), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n558), .A2(new_n559), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n232), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n526), .A2(new_n527), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n582));
  NAND2_X1  g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G71gat), .ZN(new_n585));
  INV_X1    g384(.A(G78gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT98), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT99), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n585), .B(new_n586), .C1(KEYINPUT100), .C2(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n583), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT100), .B1(new_n584), .B2(KEYINPUT9), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n581), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n563), .B1(new_n599), .B2(KEYINPUT21), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT102), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n207), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(G155gat), .B(G183gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n377), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n617), .B2(new_n406), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT103), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n621), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(KEYINPUT103), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT104), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n557), .ZN(new_n627));
  NAND3_X1  g426(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n556), .ZN(new_n629));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(KEYINPUT105), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(KEYINPUT105), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n634), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n203), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n599), .A2(new_n623), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n592), .A2(new_n598), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n624), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n648), .A2(new_n641), .A3(new_n203), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n233), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n368), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n640), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n580), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n365), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT107), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n529), .A2(new_n532), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n661), .A2(new_n458), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n529), .A2(new_n532), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n661), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n532), .B1(new_n671), .B2(new_n495), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n667), .B2(new_n666), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n673), .B2(new_n669), .ZN(G1325gat));
  AND3_X1   g473(.A1(new_n671), .A2(G15gat), .A3(new_n307), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n298), .A2(new_n299), .ZN(new_n676));
  AOI21_X1  g475(.A(G15gat), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT108), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(KEYINPUT108), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n661), .A2(new_n454), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n639), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n526), .A2(new_n527), .A3(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n510), .A2(new_n298), .A3(new_n299), .ZN(new_n687));
  INV_X1    g486(.A(new_n520), .ZN(new_n688));
  INV_X1    g487(.A(new_n521), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .A4(new_n419), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n517), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n512), .A2(new_n501), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT109), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n512), .A2(new_n501), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n684), .B1(new_n697), .B2(new_n639), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n613), .A2(new_n659), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n686), .A2(new_n698), .A3(new_n579), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n365), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n526), .A2(new_n527), .A3(new_n579), .A4(new_n699), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n365), .A3(new_n639), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(new_n543), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n703), .B2(new_n543), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT110), .B(new_n701), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1328gat));
  NOR2_X1   g510(.A1(new_n702), .A2(new_n639), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n544), .A3(new_n495), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n700), .B2(new_n458), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  NAND2_X1  g515(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n307), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n676), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n702), .A2(new_n719), .A3(new_n639), .ZN(new_n720));
  OAI221_X1 g519(.A(new_n717), .B1(new_n700), .B2(new_n718), .C1(new_n720), .C2(G43gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n721), .B(new_n722), .Z(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n700), .B2(new_n454), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n712), .A2(new_n438), .A3(new_n510), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n728), .B(new_n729), .Z(G1331gat));
  NOR2_X1   g529(.A1(new_n697), .A2(new_n579), .ZN(new_n731));
  INV_X1    g530(.A(new_n659), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n640), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n365), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n734), .A2(new_n458), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g542(.A1(new_n735), .A2(G71gat), .A3(new_n307), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n585), .B1(new_n734), .B2(new_n719), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT113), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g550(.A1(new_n734), .A2(new_n454), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n586), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n613), .A2(new_n579), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n686), .A2(new_n698), .A3(new_n659), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n365), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT114), .B1(new_n697), .B2(new_n639), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n512), .A2(new_n501), .A3(new_n695), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n695), .B1(new_n512), .B2(new_n501), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n523), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n761), .A3(new_n638), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n757), .A2(new_n762), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT115), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n763), .B2(new_n764), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n617), .B(new_n659), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n756), .B1(new_n770), .B2(new_n365), .ZN(G1336gat));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n766), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n769), .B1(new_n773), .B2(new_n768), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n732), .A2(G92gat), .A3(new_n458), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n755), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n406), .B1(new_n778), .B2(new_n495), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT116), .B(new_n775), .C1(new_n767), .C2(new_n769), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n776), .B1(new_n765), .B2(new_n766), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  XNOR2_X1  g585(.A(KEYINPUT118), .B(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n659), .A2(new_n676), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n307), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n755), .A2(new_n789), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n774), .A2(new_n788), .B1(new_n790), .B2(new_n787), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n755), .B2(new_n454), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n732), .A2(G106gat), .A3(new_n454), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n793), .C1(new_n774), .C2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n773), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n793), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(KEYINPUT53), .ZN(new_n800));
  AOI211_X1 g599(.A(KEYINPUT119), .B(new_n792), .C1(new_n798), .C2(new_n793), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(G1339gat));
  INV_X1    g601(.A(new_n579), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n660), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n652), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n650), .A2(new_n642), .A3(new_n651), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n656), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n652), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n813), .A2(new_n579), .A3(new_n657), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n558), .A2(new_n559), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n564), .A2(new_n565), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n573), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n577), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n659), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n639), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n613), .ZN(new_n822));
  AND4_X1   g621(.A1(new_n657), .A2(new_n813), .A3(new_n819), .A4(new_n814), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n821), .B(new_n822), .C1(new_n639), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n687), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n495), .A2(new_n365), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n579), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G113gat), .ZN(G1340gat));
  INV_X1    g629(.A(new_n828), .ZN(new_n831));
  OAI21_X1  g630(.A(G120gat), .B1(new_n831), .B2(new_n732), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n659), .A2(new_n214), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT120), .Z(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n831), .B2(new_n834), .ZN(G1341gat));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n613), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(G127gat), .ZN(G1342gat));
  OAI21_X1  g636(.A(G134gat), .B1(new_n831), .B2(new_n639), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n365), .B1(new_n804), .B2(new_n824), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n638), .A2(new_n458), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT121), .Z(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n839), .A2(new_n205), .A3(new_n687), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT56), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n838), .A2(new_n844), .ZN(G1343gat));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n825), .B2(new_n510), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT57), .B(new_n454), .C1(new_n804), .C2(new_n824), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n789), .A3(new_n579), .A4(new_n827), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n803), .A2(G141gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n307), .A2(new_n454), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n825), .A2(new_n736), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n495), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n851), .A2(G141gat), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT122), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n858), .A3(new_n853), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n495), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n852), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n846), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n825), .A2(new_n510), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n825), .A2(new_n847), .A3(new_n510), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(new_n789), .A3(new_n827), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n322), .B1(new_n867), .B2(new_n579), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n846), .A2(new_n856), .B1(new_n862), .B2(new_n868), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n860), .A2(new_n320), .A3(new_n659), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n789), .A3(new_n659), .A4(new_n827), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(G148gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n871), .B2(G148gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1345gat));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  AOI21_X1  g676(.A(G155gat), .B1(new_n860), .B2(new_n613), .ZN(new_n878));
  INV_X1    g677(.A(G155gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n866), .A2(new_n879), .A3(new_n822), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n857), .A2(new_n859), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n458), .A3(new_n613), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n879), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n822), .A2(new_n879), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT123), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n866), .B2(new_n639), .ZN(new_n889));
  INV_X1    g688(.A(G162gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n882), .A2(new_n890), .A3(new_n842), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1347gat));
  AOI21_X1  g691(.A(new_n736), .B1(new_n804), .B2(new_n824), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n687), .A2(KEYINPUT124), .A3(new_n495), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  INV_X1    g694(.A(new_n687), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n458), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n232), .A3(new_n579), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n893), .A2(new_n687), .A3(new_n495), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n803), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1348gat));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n233), .A3(new_n659), .ZN(new_n903));
  OAI21_X1  g702(.A(G176gat), .B1(new_n900), .B2(new_n732), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n905), .B(new_n906), .ZN(G1349gat));
  NAND4_X1  g706(.A1(new_n898), .A2(KEYINPUT126), .A3(new_n254), .A4(new_n613), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n254), .A3(new_n894), .A4(new_n897), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n822), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G183gat), .B1(new_n900), .B2(new_n822), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n900), .B2(new_n639), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n255), .A3(new_n638), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n458), .A2(new_n736), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n850), .A2(new_n789), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n803), .ZN(new_n925));
  AND4_X1   g724(.A1(new_n365), .A2(new_n825), .A3(new_n495), .A4(new_n853), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n367), .A3(new_n579), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n368), .A3(new_n659), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT62), .Z(new_n930));
  OAI21_X1  g729(.A(G204gat), .B1(new_n924), .B2(new_n732), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1353gat));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n377), .A3(new_n613), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n850), .A2(new_n789), .A3(new_n613), .A4(new_n923), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  NOR3_X1   g737(.A1(new_n924), .A2(new_n378), .A3(new_n639), .ZN(new_n939));
  AOI21_X1  g738(.A(G218gat), .B1(new_n926), .B2(new_n638), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1355gat));
endmodule


