

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n413), .B(n412), .ZN(n414) );
  NOR2_X1 U324 ( .A1(n532), .A2(n475), .ZN(n566) );
  XNOR2_X1 U325 ( .A(KEYINPUT107), .B(KEYINPUT38), .ZN(n451) );
  XOR2_X1 U326 ( .A(n324), .B(n323), .Z(n523) );
  AND2_X1 U327 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U328 ( .A(G134GAT), .B(G106GAT), .Z(n292) );
  XNOR2_X1 U329 ( .A(G99GAT), .B(G85GAT), .ZN(n403) );
  XNOR2_X1 U330 ( .A(n462), .B(KEYINPUT45), .ZN(n463) );
  XNOR2_X1 U331 ( .A(n398), .B(n291), .ZN(n318) );
  XNOR2_X1 U332 ( .A(n402), .B(n292), .ZN(n407) );
  INV_X1 U333 ( .A(KEYINPUT37), .ZN(n412) );
  XNOR2_X1 U334 ( .A(n318), .B(n388), .ZN(n319) );
  XNOR2_X1 U335 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U336 ( .A(KEYINPUT36), .B(n565), .Z(n583) );
  NOR2_X1 U337 ( .A1(n471), .A2(n520), .ZN(n570) );
  XNOR2_X1 U338 ( .A(n415), .B(n414), .ZN(n519) );
  XOR2_X1 U339 ( .A(n433), .B(n410), .Z(n565) );
  XNOR2_X1 U340 ( .A(n452), .B(n451), .ZN(n504) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U342 ( .A(n453), .B(G43GAT), .ZN(n454) );
  XNOR2_X1 U343 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G190GAT), .B(G99GAT), .Z(n294) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n297) );
  XOR2_X1 U348 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n296) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n320) );
  XOR2_X1 U351 ( .A(n297), .B(n320), .Z(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT64), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(KEYINPUT85), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U355 ( .A(G71GAT), .B(G176GAT), .Z(n301) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT0), .B(G120GAT), .Z(n307) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U363 ( .A(G134GAT), .B(KEYINPUT84), .Z(n308) );
  XOR2_X1 U364 ( .A(n309), .B(n308), .Z(n360) );
  XOR2_X1 U365 ( .A(n310), .B(n360), .Z(n532) );
  XOR2_X1 U366 ( .A(KEYINPUT21), .B(G218GAT), .Z(n312) );
  XNOR2_X1 U367 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(G197GAT), .B(n313), .Z(n329) );
  XOR2_X1 U370 ( .A(G92GAT), .B(G64GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(G204GAT), .B(KEYINPUT76), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U373 ( .A(G176GAT), .B(n316), .Z(n438) );
  XNOR2_X1 U374 ( .A(n329), .B(n438), .ZN(n324) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XNOR2_X1 U376 ( .A(G8GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n317), .B(KEYINPUT80), .ZN(n388) );
  XOR2_X1 U378 ( .A(n319), .B(KEYINPUT94), .Z(n322) );
  XNOR2_X1 U379 ( .A(n320), .B(KEYINPUT93), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  INV_X1 U381 ( .A(n523), .ZN(n468) );
  NOR2_X1 U382 ( .A1(n532), .A2(n468), .ZN(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT97), .B(n325), .ZN(n340) );
  XOR2_X1 U384 ( .A(KEYINPUT22), .B(G204GAT), .Z(n327) );
  XOR2_X1 U385 ( .A(G141GAT), .B(G22GAT), .Z(n428) );
  XOR2_X1 U386 ( .A(G50GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U387 ( .A(n428), .B(n399), .ZN(n326) );
  XOR2_X1 U388 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n331) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G78GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n332), .B(G148GAT), .ZN(n444) );
  XNOR2_X1 U394 ( .A(n333), .B(n444), .ZN(n335) );
  XNOR2_X1 U395 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U397 ( .A(KEYINPUT3), .B(KEYINPUT87), .Z(n337) );
  XNOR2_X1 U398 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(KEYINPUT2), .B(n338), .Z(n352) );
  XNOR2_X1 U401 ( .A(n339), .B(n352), .ZN(n472) );
  NAND2_X1 U402 ( .A1(n340), .A2(n472), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(KEYINPUT25), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n523), .B(KEYINPUT27), .ZN(n370) );
  INV_X1 U405 ( .A(n532), .ZN(n525) );
  NOR2_X1 U406 ( .A1(n472), .A2(n525), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n342), .B(KEYINPUT26), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n343), .B(KEYINPUT96), .ZN(n569) );
  AND2_X1 U409 ( .A1(n370), .A2(n569), .ZN(n344) );
  NOR2_X1 U410 ( .A1(n345), .A2(n344), .ZN(n367) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n347) );
  XNOR2_X1 U412 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U414 ( .A(G57GAT), .B(n348), .Z(n350) );
  NAND2_X1 U415 ( .A1(G225GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U417 ( .A(n351), .B(KEYINPUT1), .Z(n355) );
  INV_X1 U418 ( .A(n352), .ZN(n353) );
  XOR2_X1 U419 ( .A(G1GAT), .B(n353), .Z(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U421 ( .A(G85GAT), .B(G162GAT), .Z(n357) );
  XNOR2_X1 U422 ( .A(G29GAT), .B(G141GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n366) );
  INV_X1 U425 ( .A(n360), .ZN(n364) );
  XOR2_X1 U426 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n362) );
  XNOR2_X1 U427 ( .A(G148GAT), .B(KEYINPUT4), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U429 ( .A(n364), .B(n363), .Z(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n520) );
  NOR2_X1 U431 ( .A1(n367), .A2(n520), .ZN(n369) );
  INV_X1 U432 ( .A(KEYINPUT98), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n374) );
  NAND2_X1 U434 ( .A1(n520), .A2(n370), .ZN(n548) );
  XOR2_X1 U435 ( .A(n472), .B(KEYINPUT66), .Z(n371) );
  XNOR2_X1 U436 ( .A(KEYINPUT28), .B(n371), .ZN(n527) );
  NOR2_X1 U437 ( .A1(n548), .A2(n527), .ZN(n534) );
  XOR2_X1 U438 ( .A(n534), .B(KEYINPUT95), .Z(n372) );
  NAND2_X1 U439 ( .A1(n532), .A2(n372), .ZN(n373) );
  NAND2_X1 U440 ( .A1(n374), .A2(n373), .ZN(n484) );
  XOR2_X1 U441 ( .A(G15GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U442 ( .A(G78GAT), .B(G211GAT), .Z(n376) );
  XNOR2_X1 U443 ( .A(G22GAT), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U445 ( .A(n424), .B(n377), .Z(n379) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n392) );
  XOR2_X1 U448 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n381) );
  XNOR2_X1 U449 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U451 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n383) );
  XNOR2_X1 U452 ( .A(G127GAT), .B(G64GAT), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U454 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U455 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n387) );
  XNOR2_X1 U456 ( .A(G71GAT), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n439) );
  XNOR2_X1 U458 ( .A(n388), .B(n439), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n482) );
  INV_X1 U461 ( .A(n482), .ZN(n579) );
  XOR2_X1 U462 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n394) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(G29GAT), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U465 ( .A(KEYINPUT7), .B(n395), .ZN(n433) );
  XOR2_X1 U466 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n397) );
  XNOR2_X1 U467 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n396) );
  XNOR2_X1 U468 ( .A(n397), .B(n396), .ZN(n409) );
  XOR2_X1 U469 ( .A(KEYINPUT9), .B(n398), .Z(n401) );
  XNOR2_X1 U470 ( .A(G218GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(KEYINPUT75), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n442), .B(KEYINPUT11), .ZN(n405) );
  AND2_X1 U474 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U476 ( .A(n409), .B(n408), .Z(n410) );
  NOR2_X1 U477 ( .A1(n579), .A2(n583), .ZN(n411) );
  AND2_X1 U478 ( .A1(n484), .A2(n411), .ZN(n415) );
  INV_X1 U479 ( .A(KEYINPUT106), .ZN(n413) );
  INV_X1 U480 ( .A(n519), .ZN(n450) );
  XOR2_X1 U481 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n432) );
  XOR2_X1 U484 ( .A(G197GAT), .B(G36GAT), .Z(n419) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(G50GAT), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U487 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n421) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(G8GAT), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U490 ( .A(n423), .B(n422), .Z(n430) );
  XOR2_X1 U491 ( .A(n424), .B(KEYINPUT72), .Z(n426) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n507) );
  INV_X1 U498 ( .A(n507), .ZN(n571) );
  XOR2_X1 U499 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n436) );
  XNOR2_X1 U500 ( .A(KEYINPUT77), .B(KEYINPUT31), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n448) );
  XOR2_X1 U503 ( .A(n439), .B(KEYINPUT32), .Z(n441) );
  NAND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U506 ( .A(n443), .B(n442), .Z(n446) );
  XNOR2_X1 U507 ( .A(G120GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n576) );
  NAND2_X1 U510 ( .A1(n571), .A2(n576), .ZN(n449) );
  XOR2_X1 U511 ( .A(KEYINPUT78), .B(n449), .Z(n488) );
  NAND2_X1 U512 ( .A1(n450), .A2(n488), .ZN(n452) );
  NAND2_X1 U513 ( .A1(n504), .A2(n525), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT55), .B(KEYINPUT124), .ZN(n474) );
  INV_X1 U516 ( .A(KEYINPUT54), .ZN(n470) );
  INV_X1 U517 ( .A(n565), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n457) );
  XNOR2_X1 U519 ( .A(n576), .B(KEYINPUT41), .ZN(n555) );
  NAND2_X1 U520 ( .A1(n555), .A2(n571), .ZN(n456) );
  XNOR2_X1 U521 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U522 ( .A1(n579), .A2(n458), .ZN(n459) );
  NAND2_X1 U523 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n583), .A2(n482), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n463), .A2(n576), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n571), .A2(n464), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT48), .B(n467), .ZN(n551) );
  NOR2_X1 U530 ( .A1(n468), .A2(n551), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n570), .A2(n472), .ZN(n473) );
  XOR2_X1 U533 ( .A(n474), .B(n473), .Z(n475) );
  XOR2_X1 U534 ( .A(KEYINPUT111), .B(n555), .Z(n537) );
  NAND2_X1 U535 ( .A1(n566), .A2(n537), .ZN(n479) );
  XOR2_X1 U536 ( .A(G176GAT), .B(KEYINPUT57), .Z(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT125), .B(KEYINPUT56), .Z(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n491) );
  NOR2_X1 U541 ( .A1(n565), .A2(n482), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n483), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n486) );
  XOR2_X1 U544 ( .A(n486), .B(KEYINPUT99), .Z(n508) );
  INV_X1 U545 ( .A(n508), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(n489), .Z(n497) );
  NAND2_X1 U548 ( .A1(n520), .A2(n497), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(G8GAT), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U551 ( .A1(n497), .A2(n523), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U554 ( .A1(n497), .A2(n525), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT105), .Z(n499) );
  NAND2_X1 U558 ( .A1(n497), .A2(n527), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U561 ( .A1(n520), .A2(n504), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n504), .A2(n523), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT108), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n527), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n510) );
  NAND2_X1 U570 ( .A1(n507), .A2(n537), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n508), .A2(n518), .ZN(n514) );
  NAND2_X1 U572 ( .A1(n514), .A2(n520), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  NAND2_X1 U575 ( .A1(n523), .A2(n514), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n525), .A2(n514), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n516) );
  NAND2_X1 U580 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n520), .A2(n528), .ZN(n521) );
  XNOR2_X1 U585 ( .A(KEYINPUT114), .B(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n528), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n528), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n551), .A2(n532), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(KEYINPUT117), .B(n535), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n571), .A2(n545), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT118), .Z(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n543) );
  NAND2_X1 U606 ( .A1(n545), .A2(n579), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n544), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U610 ( .A1(n545), .A2(n565), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  INV_X1 U612 ( .A(n548), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n549), .A2(n569), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n561) );
  AND2_X1 U615 ( .A1(n571), .A2(n561), .ZN(n552) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n559) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U621 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n579), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n566), .A2(n571), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n579), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n571), .A2(n580), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  OR2_X1 U643 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

