

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  INV_X1 U324 ( .A(n576), .ZN(n493) );
  XOR2_X1 U325 ( .A(G113GAT), .B(KEYINPUT0), .Z(n347) );
  XNOR2_X1 U326 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X1 U327 ( .A(n353), .ZN(n354) );
  OR2_X1 U328 ( .A1(n483), .A2(n478), .ZN(n479) );
  XNOR2_X1 U329 ( .A(n309), .B(n308), .ZN(n589) );
  XOR2_X1 U330 ( .A(KEYINPUT38), .B(n452), .Z(n514) );
  XNOR2_X1 U331 ( .A(n373), .B(n372), .ZN(n375) );
  XNOR2_X1 U332 ( .A(n371), .B(n370), .ZN(n372) );
  AND2_X1 U333 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U334 ( .A(n300), .B(n299), .Z(n293) );
  XOR2_X1 U335 ( .A(n438), .B(n329), .Z(n294) );
  INV_X1 U336 ( .A(KEYINPUT95), .ZN(n376) );
  XNOR2_X1 U337 ( .A(n377), .B(n376), .ZN(n378) );
  INV_X1 U338 ( .A(KEYINPUT25), .ZN(n379) );
  XNOR2_X1 U339 ( .A(n380), .B(n379), .ZN(n384) );
  NOR2_X1 U340 ( .A1(n465), .A2(n586), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n392), .B(KEYINPUT9), .ZN(n393) );
  XNOR2_X1 U342 ( .A(n473), .B(KEYINPUT120), .ZN(n474) );
  XNOR2_X1 U343 ( .A(n394), .B(n393), .ZN(n401) );
  XNOR2_X1 U344 ( .A(n301), .B(n293), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n409), .B(n292), .ZN(n365) );
  XNOR2_X1 U346 ( .A(n475), .B(n474), .ZN(n483) );
  XNOR2_X1 U347 ( .A(n401), .B(n447), .ZN(n404) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n365), .B(n364), .ZN(n366) );
  NOR2_X1 U350 ( .A1(n531), .A2(n483), .ZN(n484) );
  INV_X1 U351 ( .A(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U352 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U353 ( .A(n435), .B(n410), .ZN(n411) );
  OR2_X1 U354 ( .A1(n529), .A2(n501), .ZN(n452) );
  XNOR2_X1 U355 ( .A(n485), .B(KEYINPUT126), .ZN(n590) );
  XNOR2_X1 U356 ( .A(n412), .B(n411), .ZN(n572) );
  XNOR2_X1 U357 ( .A(n363), .B(n374), .ZN(n542) );
  XNOR2_X1 U358 ( .A(KEYINPUT62), .B(G218GAT), .ZN(n487) );
  XNOR2_X1 U359 ( .A(n494), .B(G190GAT), .ZN(n495) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U361 ( .A(n488), .B(n487), .ZN(G1355GAT) );
  XNOR2_X1 U362 ( .A(n496), .B(n495), .ZN(G1351GAT) );
  XNOR2_X1 U363 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U364 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n296) );
  XNOR2_X1 U365 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n295) );
  XNOR2_X1 U366 ( .A(n296), .B(n295), .ZN(n309) );
  XNOR2_X1 U367 ( .A(G57GAT), .B(G64GAT), .ZN(n297) );
  XNOR2_X1 U368 ( .A(n297), .B(KEYINPUT13), .ZN(n438) );
  XOR2_X1 U369 ( .A(G22GAT), .B(G155GAT), .Z(n329) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U371 ( .A(n294), .B(n298), .ZN(n303) );
  XOR2_X1 U372 ( .A(G1GAT), .B(KEYINPUT71), .Z(n422) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n353) );
  XNOR2_X1 U374 ( .A(n422), .B(n353), .ZN(n301) );
  XOR2_X1 U375 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n300) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G78GAT), .ZN(n299) );
  XOR2_X1 U377 ( .A(n304), .B(KEYINPUT81), .Z(n307) );
  XNOR2_X1 U378 ( .A(G8GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U379 ( .A(n305), .B(G211GAT), .ZN(n364) );
  XNOR2_X1 U380 ( .A(n364), .B(KEYINPUT80), .ZN(n306) );
  XNOR2_X1 U381 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U382 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n311) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n310) );
  XNOR2_X1 U384 ( .A(n311), .B(n310), .ZN(n330) );
  XOR2_X1 U385 ( .A(n330), .B(KEYINPUT5), .Z(n313) );
  NAND2_X1 U386 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U387 ( .A(n313), .B(n312), .ZN(n328) );
  XOR2_X1 U388 ( .A(G57GAT), .B(G120GAT), .Z(n315) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U390 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U391 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n317) );
  XNOR2_X1 U392 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n316) );
  XNOR2_X1 U393 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U394 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U395 ( .A(G155GAT), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U396 ( .A(G134GAT), .B(G148GAT), .ZN(n320) );
  XNOR2_X1 U397 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U398 ( .A(n322), .B(G85GAT), .Z(n324) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(n347), .ZN(n323) );
  XNOR2_X1 U400 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U401 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U402 ( .A(n328), .B(n327), .ZN(n531) );
  XOR2_X1 U403 ( .A(n330), .B(n329), .Z(n332) );
  NAND2_X1 U404 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U405 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U406 ( .A(n333), .B(G211GAT), .Z(n337) );
  XOR2_X1 U407 ( .A(G162GAT), .B(KEYINPUT76), .Z(n335) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U409 ( .A(n335), .B(n334), .ZN(n402) );
  XNOR2_X1 U410 ( .A(n402), .B(KEYINPUT22), .ZN(n336) );
  XNOR2_X1 U411 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n339) );
  XNOR2_X1 U413 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n338) );
  XNOR2_X1 U414 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U415 ( .A(n341), .B(n340), .Z(n346) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n342) );
  XNOR2_X1 U417 ( .A(n342), .B(KEYINPUT21), .ZN(n367) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G148GAT), .Z(n344) );
  XNOR2_X1 U419 ( .A(KEYINPUT73), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U420 ( .A(n344), .B(n343), .ZN(n439) );
  XNOR2_X1 U421 ( .A(n367), .B(n439), .ZN(n345) );
  XNOR2_X1 U422 ( .A(n346), .B(n345), .ZN(n476) );
  XOR2_X1 U423 ( .A(G120GAT), .B(G71GAT), .Z(n443) );
  XOR2_X1 U424 ( .A(n443), .B(n347), .Z(n349) );
  NAND2_X1 U425 ( .A1(G227GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U426 ( .A(n349), .B(n348), .ZN(n357) );
  XOR2_X1 U427 ( .A(G183GAT), .B(KEYINPUT84), .Z(n351) );
  XNOR2_X1 U428 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n350) );
  XNOR2_X1 U429 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U430 ( .A(G43GAT), .B(G134GAT), .Z(n394) );
  XNOR2_X1 U431 ( .A(n352), .B(n394), .ZN(n355) );
  XNOR2_X1 U432 ( .A(G190GAT), .B(G99GAT), .ZN(n358) );
  XNOR2_X1 U433 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U434 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n361) );
  XNOR2_X1 U435 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n360) );
  XNOR2_X1 U436 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(n362), .ZN(n374) );
  XOR2_X1 U438 ( .A(G36GAT), .B(G190GAT), .Z(n409) );
  XOR2_X1 U439 ( .A(n366), .B(KEYINPUT91), .Z(n373) );
  XNOR2_X1 U440 ( .A(n367), .B(G64GAT), .ZN(n371) );
  XOR2_X1 U441 ( .A(KEYINPUT92), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U442 ( .A(G204GAT), .B(G218GAT), .ZN(n368) );
  XNOR2_X1 U443 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n533) );
  NAND2_X1 U445 ( .A1(n542), .A2(n533), .ZN(n377) );
  NAND2_X1 U446 ( .A1(n476), .A2(n378), .ZN(n380) );
  XNOR2_X1 U447 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n382) );
  NOR2_X1 U448 ( .A1(n542), .A2(n476), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n558) );
  XNOR2_X1 U450 ( .A(KEYINPUT27), .B(n533), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n558), .A2(n387), .ZN(n383) );
  NAND2_X1 U452 ( .A1(n384), .A2(n383), .ZN(n385) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(n385), .Z(n386) );
  NOR2_X1 U454 ( .A1(n531), .A2(n386), .ZN(n391) );
  NAND2_X1 U455 ( .A1(n531), .A2(n387), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n388), .B(KEYINPUT93), .ZN(n557) );
  XNOR2_X1 U457 ( .A(n476), .B(KEYINPUT28), .ZN(n509) );
  NAND2_X1 U458 ( .A1(n557), .A2(n509), .ZN(n544) );
  XNOR2_X1 U459 ( .A(KEYINPUT86), .B(n542), .ZN(n389) );
  NOR2_X1 U460 ( .A1(n544), .A2(n389), .ZN(n390) );
  NOR2_X1 U461 ( .A1(n391), .A2(n390), .ZN(n499) );
  INV_X1 U462 ( .A(KEYINPUT78), .ZN(n413) );
  AND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  INV_X1 U464 ( .A(G85GAT), .ZN(n395) );
  NAND2_X1 U465 ( .A1(G92GAT), .A2(n395), .ZN(n398) );
  INV_X1 U466 ( .A(G92GAT), .ZN(n396) );
  NAND2_X1 U467 ( .A1(n396), .A2(G85GAT), .ZN(n397) );
  NAND2_X1 U468 ( .A1(n398), .A2(n397), .ZN(n400) );
  XNOR2_X1 U469 ( .A(G99GAT), .B(G106GAT), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n447) );
  XOR2_X1 U471 ( .A(n402), .B(KEYINPUT77), .Z(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n405), .B(KEYINPUT10), .ZN(n412) );
  XOR2_X1 U474 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n407) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U477 ( .A(KEYINPUT7), .B(n408), .Z(n435) );
  XOR2_X1 U478 ( .A(n409), .B(KEYINPUT11), .Z(n410) );
  XNOR2_X1 U479 ( .A(n413), .B(n572), .ZN(n492) );
  XOR2_X1 U480 ( .A(KEYINPUT36), .B(n492), .Z(n486) );
  NOR2_X1 U481 ( .A1(n499), .A2(n486), .ZN(n414) );
  NAND2_X1 U482 ( .A1(n589), .A2(n414), .ZN(n415) );
  XOR2_X1 U483 ( .A(n415), .B(KEYINPUT37), .Z(n529) );
  XOR2_X1 U484 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n417) );
  XNOR2_X1 U485 ( .A(G15GAT), .B(G8GAT), .ZN(n416) );
  XNOR2_X1 U486 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U487 ( .A(KEYINPUT66), .B(KEYINPUT72), .Z(n419) );
  XNOR2_X1 U488 ( .A(KEYINPUT65), .B(KEYINPUT29), .ZN(n418) );
  XNOR2_X1 U489 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U490 ( .A(n421), .B(n420), .Z(n427) );
  XOR2_X1 U491 ( .A(KEYINPUT30), .B(n422), .Z(n424) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U494 ( .A(KEYINPUT64), .B(n425), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U496 ( .A(G197GAT), .B(G36GAT), .Z(n429) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(G43GAT), .ZN(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U499 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U500 ( .A(G113GAT), .B(G22GAT), .Z(n433) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G141GAT), .ZN(n432) );
  XNOR2_X1 U502 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U504 ( .A(n437), .B(n436), .ZN(n581) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n451) );
  XOR2_X1 U506 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n441) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n440) );
  XNOR2_X1 U508 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U509 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U510 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U511 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U512 ( .A(n446), .B(KEYINPUT32), .Z(n449) );
  XNOR2_X1 U513 ( .A(n447), .B(KEYINPUT74), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U515 ( .A(n451), .B(n450), .ZN(n586) );
  OR2_X1 U516 ( .A1(n581), .A2(n586), .ZN(n501) );
  NAND2_X1 U517 ( .A1(n514), .A2(n542), .ZN(n454) );
  NAND2_X1 U518 ( .A1(n514), .A2(n531), .ZN(n457) );
  XOR2_X1 U519 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n455) );
  XNOR2_X1 U520 ( .A(n455), .B(G29GAT), .ZN(n456) );
  XNOR2_X1 U521 ( .A(n457), .B(n456), .ZN(G1328GAT) );
  XOR2_X1 U522 ( .A(KEYINPUT111), .B(KEYINPUT47), .Z(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT109), .B(n589), .ZN(n549) );
  XNOR2_X1 U524 ( .A(KEYINPUT41), .B(n586), .ZN(n575) );
  NOR2_X1 U525 ( .A1(n581), .A2(n575), .ZN(n458) );
  XNOR2_X1 U526 ( .A(KEYINPUT46), .B(n458), .ZN(n459) );
  XNOR2_X1 U527 ( .A(KEYINPUT110), .B(n459), .ZN(n460) );
  NOR2_X1 U528 ( .A1(n549), .A2(n460), .ZN(n461) );
  NAND2_X1 U529 ( .A1(n461), .A2(n572), .ZN(n462) );
  XNOR2_X1 U530 ( .A(n463), .B(n462), .ZN(n470) );
  INV_X1 U531 ( .A(n581), .ZN(n561) );
  NOR2_X1 U532 ( .A1(n589), .A2(n486), .ZN(n464) );
  XOR2_X1 U533 ( .A(KEYINPUT45), .B(n464), .Z(n465) );
  XNOR2_X1 U534 ( .A(n466), .B(KEYINPUT112), .ZN(n467) );
  AND2_X1 U535 ( .A1(n581), .A2(n467), .ZN(n468) );
  XOR2_X1 U536 ( .A(KEYINPUT113), .B(n468), .Z(n469) );
  NOR2_X2 U537 ( .A1(n470), .A2(n469), .ZN(n472) );
  XNOR2_X2 U538 ( .A(n472), .B(n471), .ZN(n560) );
  NAND2_X1 U539 ( .A1(n560), .A2(n533), .ZN(n475) );
  XOR2_X1 U540 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n473) );
  INV_X1 U541 ( .A(n531), .ZN(n477) );
  NAND2_X1 U542 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(KEYINPUT55), .ZN(n480) );
  NAND2_X1 U544 ( .A1(n480), .A2(n542), .ZN(n576) );
  NAND2_X1 U545 ( .A1(n493), .A2(n549), .ZN(n482) );
  XNOR2_X1 U546 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n481) );
  XNOR2_X1 U547 ( .A(n482), .B(n481), .ZN(G1350GAT) );
  NAND2_X1 U548 ( .A1(n558), .A2(n484), .ZN(n485) );
  OR2_X1 U549 ( .A1(n590), .A2(n486), .ZN(n488) );
  NOR2_X1 U550 ( .A1(n581), .A2(n576), .ZN(n491) );
  INV_X1 U551 ( .A(G169GAT), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT122), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1348GAT) );
  AND2_X1 U554 ( .A1(n493), .A2(n492), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n589), .A2(n492), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT16), .B(n497), .Z(n498) );
  NOR2_X1 U558 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(n500), .ZN(n517) );
  NOR2_X1 U560 ( .A1(n501), .A2(n517), .ZN(n510) );
  NAND2_X1 U561 ( .A1(n531), .A2(n510), .ZN(n504) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT98), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n533), .A2(n510), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U568 ( .A1(n510), .A2(n542), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U570 ( .A(G15GAT), .B(n508), .Z(G1326GAT) );
  INV_X1 U571 ( .A(n509), .ZN(n538) );
  NAND2_X1 U572 ( .A1(n510), .A2(n538), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U574 ( .A(G36GAT), .B(KEYINPUT101), .Z(n513) );
  NAND2_X1 U575 ( .A1(n514), .A2(n533), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n538), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n519) );
  INV_X1 U580 ( .A(n575), .ZN(n563) );
  NAND2_X1 U581 ( .A1(n563), .A2(n581), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(KEYINPUT102), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n530), .A2(n517), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n525), .A2(n531), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n533), .A2(n525), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT104), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G64GAT), .B(n522), .ZN(G1333GAT) );
  XOR2_X1 U590 ( .A(G71GAT), .B(KEYINPUT105), .Z(n524) );
  NAND2_X1 U591 ( .A1(n525), .A2(n542), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U594 ( .A1(n525), .A2(n538), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n539), .A2(n531), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  XOR2_X1 U600 ( .A(G92GAT), .B(KEYINPUT107), .Z(n535) );
  NAND2_X1 U601 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1337GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n542), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT108), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G99GAT), .B(n537), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n540), .B(KEYINPUT44), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n560), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n561), .A2(n553), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U614 ( .A1(n553), .A2(n563), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n551) );
  NAND2_X1 U618 ( .A1(n553), .A2(n549), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n555) );
  NAND2_X1 U622 ( .A1(n553), .A2(n492), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G134GAT), .B(n556), .ZN(G1343GAT) );
  AND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n571) );
  INV_X1 U627 ( .A(n571), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(G148GAT), .B(KEYINPUT53), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1345GAT) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(KEYINPUT118), .ZN(n570) );
  OR2_X1 U636 ( .A1(n589), .A2(n571), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1346GAT) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1347GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n578) );
  XNOR2_X1 U643 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1349GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n590), .ZN(n584) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  INV_X1 U651 ( .A(n590), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n591), .Z(G1354GAT) );
endmodule

