//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n207), .B2(KEYINPUT87), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT87), .B2(new_n207), .ZN(new_n209));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n206), .A2(KEYINPUT88), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(KEYINPUT88), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n203), .A2(new_n210), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n220), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n211), .B2(new_n217), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n219), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n218), .A2(new_n226), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n226), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n226), .A3(KEYINPUT89), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n230), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n242), .A3(new_n248), .A4(new_n235), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT78), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(G113gat), .B2(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n260), .A2(G127gat), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n266), .A2(new_n268), .B1(KEYINPUT67), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n259), .B2(new_n261), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n258), .A2(G134gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n275), .A3(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n268), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT68), .B(G113gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n265), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n272), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n268), .B1(new_n285), .B2(G120gat), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n274), .A4(new_n276), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n271), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(KEYINPUT2), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n293), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n297), .B(new_n296), .C1(new_n303), .C2(KEYINPUT2), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n257), .B1(new_n288), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n288), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n281), .A2(new_n287), .ZN(new_n316));
  INV_X1    g115(.A(new_n271), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n313), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n311), .A3(new_n313), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n254), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n323));
  AOI211_X1 g122(.A(new_n271), .B(new_n312), .C1(new_n281), .C2(new_n287), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n256), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT80), .B(new_n256), .C1(new_n323), .C2(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n257), .A2(new_n254), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n288), .A2(new_n308), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n331), .B(new_n332), .C1(new_n319), .C2(new_n320), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G1gat), .B(G29gat), .Z(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n340), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n330), .A2(new_n342), .A3(new_n334), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n333), .B1(new_n322), .B2(new_n329), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n342), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT22), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(KEYINPUT74), .B1(G211gat), .B2(G218gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(KEYINPUT74), .B2(new_n349), .ZN(new_n351));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT76), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT75), .B1(new_n351), .B2(new_n352), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n354), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NOR4_X1   g160(.A1(new_n361), .A2(new_n357), .A3(KEYINPUT76), .A4(new_n354), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  NOR4_X1   g164(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT66), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G183gat), .ZN(new_n373));
  INV_X1    g172(.A(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT27), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(KEYINPUT64), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G183gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT27), .ZN(new_n382));
  OR3_X1    g181(.A1(new_n374), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(KEYINPUT65), .ZN(new_n384));
  NOR2_X1   g183(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT64), .B(G183gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT24), .B1(new_n374), .B2(new_n376), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT24), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n388), .A2(new_n376), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n368), .A2(KEYINPUT23), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(G169gat), .B2(G176gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n364), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT25), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(KEYINPUT25), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(new_n391), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n387), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n387), .A2(new_n397), .A3(new_n401), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT29), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n363), .B(new_n404), .C1(new_n406), .C2(new_n403), .ZN(new_n407));
  INV_X1    g206(.A(new_n357), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT76), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n359), .A4(new_n355), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n361), .A2(new_n357), .A3(new_n354), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(new_n356), .ZN(new_n412));
  INV_X1    g211(.A(new_n404), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n402), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n416), .A3(new_n420), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n407), .A2(new_n416), .A3(new_n425), .A4(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n348), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G22gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n410), .C1(new_n411), .C2(new_n356), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n313), .B1(new_n435), .B2(new_n305), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n307), .A2(new_n414), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n412), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n433), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n353), .B(new_n354), .ZN(new_n441));
  INV_X1    g240(.A(new_n414), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n305), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n312), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n444), .A3(new_n432), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT31), .B(G50gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n439), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n439), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n431), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n439), .A2(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n446), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n439), .A2(new_n445), .A3(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n430), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n316), .A2(new_n317), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n405), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n288), .A2(new_n402), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n462), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n470), .A3(new_n460), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n472));
  AND2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT72), .ZN(new_n475));
  XNOR2_X1  g274(.A(G71gat), .B(G99gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n467), .B(new_n469), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(KEYINPUT32), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n471), .B2(new_n472), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n468), .B1(new_n461), .B2(new_n462), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n470), .B(new_n466), .C1(new_n459), .C2(new_n460), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n478), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n478), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n457), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n479), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n478), .A2(new_n480), .A3(new_n484), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT36), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n456), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT6), .B1(new_n346), .B2(new_n342), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n340), .B1(new_n346), .B2(KEYINPUT84), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n496), .B(new_n333), .C1(new_n322), .C2(new_n329), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n423), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT37), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n406), .A2(new_n403), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n413), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n502), .B2(new_n412), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n363), .B1(new_n413), .B2(new_n415), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT38), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n422), .B1(new_n500), .B2(new_n420), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n498), .A2(new_n341), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n498), .A2(new_n510), .A3(new_n341), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n417), .A2(KEYINPUT37), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT38), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n450), .A2(new_n454), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n424), .A2(KEYINPUT82), .A3(new_n426), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT82), .B1(new_n424), .B2(new_n426), .ZN(new_n519));
  INV_X1    g318(.A(new_n332), .ZN(new_n520));
  INV_X1    g319(.A(new_n320), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(new_n314), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n256), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n319), .A2(new_n320), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n257), .B1(new_n525), .B2(new_n520), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n323), .A2(new_n324), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT39), .B1(new_n527), .B2(new_n256), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n342), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT40), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n518), .A2(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n495), .A2(new_n497), .B1(new_n531), .B2(new_n529), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n493), .B1(new_n515), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n489), .A2(new_n454), .A3(new_n450), .A4(new_n490), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n427), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n517), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n498), .A2(new_n341), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n485), .A2(new_n486), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n348), .A2(new_n516), .A3(new_n548), .A4(new_n427), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT86), .B1(new_n549), .B2(KEYINPUT35), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n253), .B1(new_n539), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT91), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n560), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT7), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n567), .A2(new_n568), .B1(KEYINPUT8), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n563), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n563), .A2(new_n566), .A3(new_n572), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n559), .B1(new_n218), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n219), .A2(new_n228), .A3(new_n576), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n580), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n558), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n557), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G78gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(new_n599), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n574), .A3(new_n575), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT94), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(new_n608), .A3(new_n602), .A4(new_n604), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n604), .A2(new_n602), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n595), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n601), .A2(new_n604), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n595), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n594), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(KEYINPUT95), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n594), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n612), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G127gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n226), .B1(new_n600), .B2(new_n625), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT90), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(new_n294), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n635), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n591), .A2(new_n624), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n554), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n348), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT97), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  INV_X1    g447(.A(new_n543), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n225), .B2(new_n650), .ZN(new_n653));
  MUX2_X1   g452(.A(new_n652), .B(new_n653), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n644), .B2(new_n492), .ZN(new_n655));
  INV_X1    g454(.A(new_n548), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n644), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n644), .A2(new_n516), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n642), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(new_n624), .A3(new_n253), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n667), .B2(new_n550), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT44), .B(new_n591), .C1(new_n668), .C2(new_n538), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n515), .A2(new_n537), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n346), .A2(new_n344), .A3(new_n342), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n335), .A2(new_n340), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n494), .ZN(new_n673));
  INV_X1    g472(.A(new_n427), .ZN(new_n674));
  OAI211_X1 g473(.A(KEYINPUT101), .B(new_n455), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n492), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT101), .B1(new_n428), .B2(new_n455), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n590), .B1(new_n679), .B2(new_n553), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n663), .B(new_n669), .C1(new_n680), .C2(KEYINPUT44), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n514), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n508), .B2(KEYINPUT85), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n536), .B1(new_n685), .B2(new_n511), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n494), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n674), .B1(new_n688), .B2(new_n341), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n516), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n492), .A3(new_n675), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n591), .B1(new_n692), .B2(new_n668), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n695), .A2(KEYINPUT102), .A3(new_n663), .A4(new_n669), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n683), .A2(new_n673), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n696), .A3(new_n699), .A4(new_n673), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(G29gat), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n591), .B(new_n663), .C1(new_n668), .C2(new_n538), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n705));
  INV_X1    g504(.A(G29gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n673), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT100), .B1(new_n703), .B2(new_n707), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n702), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n711), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n712), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT104), .B1(new_n701), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n698), .A2(G29gat), .A3(new_n700), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n718), .A4(new_n715), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1328gat));
  AND2_X1   g523(.A1(new_n683), .A2(new_n696), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n543), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G36gat), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n703), .A2(G36gat), .A3(new_n649), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1329gat));
  OAI21_X1  g529(.A(G43gat), .B1(new_n681), .B2(new_n492), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n703), .A2(G43gat), .A3(new_n656), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n492), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n732), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n683), .A2(new_n455), .A3(new_n696), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n516), .A2(G50gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT105), .ZN(new_n743));
  NOR4_X1   g542(.A1(new_n743), .A2(new_n662), .A3(new_n590), .A4(new_n624), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT48), .B1(new_n554), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G50gat), .B1(new_n681), .B2(new_n516), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n554), .A2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n741), .A2(new_n745), .B1(KEYINPUT48), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT106), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n679), .A2(new_n553), .ZN(new_n751));
  INV_X1    g550(.A(new_n624), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n752), .A2(new_n591), .A3(new_n642), .A4(new_n252), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n673), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT108), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(G57gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n543), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  NAND3_X1  g561(.A1(new_n754), .A2(G71gat), .A3(new_n736), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT109), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n754), .A2(new_n548), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(G71gat), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n455), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g568(.A1(new_n695), .A2(new_n669), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n662), .A2(new_n252), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n624), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n348), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n680), .A2(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n680), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n772), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n624), .A2(new_n568), .A3(new_n673), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT111), .Z(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n774), .A2(new_n784), .ZN(G1336gat));
  NAND2_X1  g584(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n776), .B(new_n786), .Z(new_n787));
  NOR3_X1   g586(.A1(new_n752), .A2(new_n649), .A3(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n543), .A3(new_n624), .A4(new_n772), .ZN(new_n790));
  INV_X1    g589(.A(new_n567), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(KEYINPUT112), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n790), .B2(new_n791), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n788), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n773), .B2(new_n492), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n752), .A2(G99gat), .A3(new_n656), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1338gat));
  NAND4_X1  g604(.A1(new_n771), .A2(new_n455), .A3(new_n624), .A4(new_n772), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n752), .A2(G106gat), .A3(new_n516), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n787), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n806), .B2(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n781), .A2(new_n808), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n240), .A2(new_n241), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n247), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n251), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n624), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n595), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n606), .A2(new_n824), .A3(new_n610), .A4(new_n609), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n609), .A2(new_n610), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n824), .A4(new_n606), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n826), .A2(new_n829), .A3(new_n612), .A4(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n827), .B2(new_n606), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n594), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n623), .A2(new_n834), .A3(new_n252), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n830), .B2(new_n833), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n591), .B1(new_n823), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n821), .A2(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n821), .A2(KEYINPUT118), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n840), .A2(new_n589), .A3(new_n587), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n623), .A2(new_n834), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n642), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n643), .A2(new_n253), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n673), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n540), .A3(new_n543), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n279), .A3(new_n252), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n455), .B1(new_n845), .B2(new_n846), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n851), .A2(new_n673), .A3(new_n548), .A4(new_n649), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n253), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1340gat));
  NAND2_X1  g653(.A1(new_n624), .A2(new_n265), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT119), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G120gat), .B1(new_n852), .B2(new_n752), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1341gat));
  NAND3_X1  g658(.A1(new_n849), .A2(new_n258), .A3(new_n662), .ZN(new_n860));
  OAI21_X1  g659(.A(G127gat), .B1(new_n852), .B2(new_n642), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT120), .Z(G1342gat));
  NAND3_X1  g662(.A1(new_n849), .A2(new_n260), .A3(new_n591), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n852), .B2(new_n590), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n492), .A2(new_n455), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n543), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n253), .A2(G141gat), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n673), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT122), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n842), .A2(new_n836), .A3(new_n843), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n843), .A2(new_n253), .A3(new_n836), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n821), .B1(new_n618), .B2(new_n623), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n590), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n662), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n643), .A2(new_n253), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n874), .B(new_n455), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n649), .A2(new_n673), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n736), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n837), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n836), .A2(KEYINPUT121), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n835), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n591), .B1(new_n887), .B2(new_n823), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n642), .B1(new_n888), .B2(new_n844), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n516), .B1(new_n889), .B2(new_n846), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n881), .B(new_n883), .C1(new_n890), .C2(new_n874), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n253), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n872), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n836), .B(new_n884), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n877), .B1(new_n897), .B2(new_n835), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n875), .B1(new_n898), .B2(new_n591), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n880), .B1(new_n899), .B2(new_n642), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n516), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(new_n252), .A3(new_n881), .A4(new_n883), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n896), .B1(new_n902), .B2(G141gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT123), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n905), .B(new_n896), .C1(new_n902), .C2(G141gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n894), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT124), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n894), .B(new_n909), .C1(new_n904), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n912), .B(G148gat), .C1(new_n891), .C2(new_n752), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n847), .A2(KEYINPUT57), .A3(new_n455), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(KEYINPUT57), .B2(new_n890), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n752), .A2(new_n736), .A3(new_n882), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n291), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n848), .A2(new_n543), .A3(new_n869), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n291), .A3(new_n624), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n891), .B2(new_n642), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n294), .A3(new_n662), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  NOR3_X1   g723(.A1(new_n891), .A2(new_n295), .A3(new_n590), .ZN(new_n925));
  AOI21_X1  g724(.A(G162gat), .B1(new_n919), .B2(new_n591), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NAND4_X1  g726(.A1(new_n851), .A2(new_n348), .A3(new_n548), .A4(new_n543), .ZN(new_n928));
  INV_X1    g727(.A(G169gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(new_n253), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n673), .B1(new_n845), .B2(new_n846), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n649), .A2(new_n540), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  AND2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n252), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n930), .A2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n928), .A2(new_n937), .A3(new_n752), .ZN(new_n938));
  AOI21_X1  g737(.A(G176gat), .B1(new_n934), .B2(new_n624), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(G1349gat));
  NAND4_X1  g739(.A1(new_n934), .A2(new_n373), .A3(new_n375), .A4(new_n662), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n928), .A2(new_n642), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n388), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n928), .B2(new_n590), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n934), .A2(new_n376), .A3(new_n591), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1351gat));
  AND4_X1   g747(.A1(new_n455), .A2(new_n931), .A3(new_n543), .A4(new_n492), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT126), .B(G197gat), .Z(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n252), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n915), .A2(new_n348), .A3(new_n543), .A4(new_n492), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n253), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n950), .ZN(G1352gat));
  INV_X1    g753(.A(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n955), .A3(new_n624), .ZN(new_n956));
  XOR2_X1   g755(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n952), .B2(new_n752), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(G211gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n949), .A2(new_n961), .A3(new_n662), .ZN(new_n962));
  OAI21_X1  g761(.A(G211gat), .B1(new_n952), .B2(new_n642), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n952), .B2(new_n590), .ZN(new_n968));
  INV_X1    g767(.A(G218gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n969), .A3(new_n591), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1355gat));
endmodule


