//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  AND4_X1   g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .A4(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n191), .B2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G128), .B1(new_n194), .B2(new_n188), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n189), .A2(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n194), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n198), .A2(new_n205), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n202), .B1(new_n201), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G224), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n212));
  XOR2_X1   g026(.A(new_n209), .B(new_n212), .Z(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n217), .A2(new_n218), .B1(KEYINPUT2), .B2(G113), .ZN(new_n219));
  XNOR2_X1  g033(.A(G116), .B(G119), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G104), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G107), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(G104), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G101), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n227), .A2(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n226), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT79), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n229), .A2(new_n243), .A3(new_n238), .A4(new_n233), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n235), .B1(new_n234), .B2(G101), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n237), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G110), .B(G122), .ZN(new_n249));
  OAI21_X1  g063(.A(G101), .B1(new_n228), .B2(new_n225), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n238), .B1(new_n231), .B2(new_n239), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT80), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n242), .A2(new_n244), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n220), .A2(KEYINPUT5), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n257), .A2(KEYINPUT5), .A3(G119), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(new_n216), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n221), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n248), .A2(new_n249), .A3(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n213), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n249), .B(KEYINPUT8), .ZN(new_n264));
  INV_X1    g078(.A(new_n261), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n255), .A2(new_n260), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n249), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n237), .A2(new_n247), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n262), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n269), .C1(new_n270), .C2(new_n265), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n209), .B(new_n211), .Z(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n268), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n268), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  INV_X1    g095(.A(G237), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n210), .A3(G214), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(G143), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT18), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n283), .B(new_n191), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT18), .A3(G131), .ZN(new_n289));
  INV_X1    g103(.A(G140), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G125), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n201), .A2(G140), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(new_n189), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT85), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT85), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n287), .A2(new_n289), .A3(new_n294), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT72), .B1(new_n291), .B2(KEYINPUT16), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(G146), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT86), .B1(new_n288), .B2(G131), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n284), .A2(new_n307), .A3(new_n286), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n288), .A2(G131), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n306), .A2(new_n308), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n304), .A2(G146), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n288), .A2(KEYINPUT17), .A3(G131), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n305), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G113), .B(G122), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n227), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n299), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n299), .B2(new_n314), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n281), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G475), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n306), .A2(new_n310), .A3(new_n308), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n293), .B(KEYINPUT19), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n323), .B(new_n312), .C1(G146), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n299), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n316), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n317), .ZN(new_n330));
  NOR2_X1   g144(.A1(G475), .A2(G902), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n322), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT20), .B(new_n333), .C1(new_n329), .C2(new_n317), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n321), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G952), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G953), .ZN(new_n338));
  INV_X1    g152(.A(G234), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n282), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n281), .B(new_n210), .C1(G234), .C2(G237), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT21), .B(G898), .Z(new_n343));
  OAI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G478), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT15), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(KEYINPUT15), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n191), .A2(G128), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT89), .ZN(new_n352));
  INV_X1    g166(.A(G134), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n191), .A2(G128), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT88), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n353), .B1(new_n352), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT91), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n358), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n356), .ZN(new_n362));
  INV_X1    g176(.A(G122), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n363), .A2(KEYINPUT87), .A3(G116), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n363), .B2(G116), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n364), .A2(new_n365), .B1(G116), .B2(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(G116), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n224), .B1(new_n367), .B2(KEYINPUT14), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n366), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n359), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT13), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n352), .B1(new_n355), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n355), .A2(new_n371), .ZN(new_n373));
  OAI21_X1  g187(.A(G134), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n357), .A2(KEYINPUT90), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n366), .B(new_n224), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n356), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT9), .B(G234), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n380), .A2(new_n381), .A3(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n370), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n370), .B2(new_n379), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n350), .B1(new_n386), .B2(G902), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n379), .ZN(new_n388));
  INV_X1    g202(.A(new_n382), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n383), .ZN(new_n391));
  INV_X1    g205(.A(new_n350), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n281), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n336), .A2(new_n344), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n280), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT11), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n353), .B2(G137), .ZN(new_n399));
  INV_X1    g213(.A(G137), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT11), .A3(G134), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n353), .A2(G137), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n286), .A4(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n353), .A2(G137), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n400), .A2(G134), .ZN(new_n405));
  OAI21_X1  g219(.A(G131), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT66), .B1(new_n200), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G131), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n403), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n208), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n403), .A2(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT66), .ZN(new_n414));
  INV_X1    g228(.A(G128), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n190), .B1(new_n206), .B2(new_n196), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n195), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n413), .B(new_n414), .C1(new_n418), .C2(new_n193), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n408), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT30), .ZN(new_n421));
  INV_X1    g235(.A(new_n200), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n413), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n412), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n223), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n419), .A2(new_n412), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n221), .A2(new_n222), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(KEYINPUT67), .A3(new_n429), .A4(new_n408), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n408), .A2(new_n429), .A3(new_n419), .A4(new_n412), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n282), .A2(new_n210), .A3(G210), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT69), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G101), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT28), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n423), .A2(new_n412), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n223), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n223), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n434), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n443), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  INV_X1    g265(.A(new_n446), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n420), .B2(new_n223), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n420), .A2(new_n223), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n434), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(new_n457), .B2(KEYINPUT28), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n441), .A2(KEYINPUT29), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G472), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n449), .B1(new_n434), .B2(new_n447), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n442), .B1(new_n463), .B2(new_n452), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT31), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n427), .A2(new_n465), .A3(new_n441), .A4(new_n434), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n427), .A2(new_n441), .A3(new_n434), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT31), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G472), .A2(G902), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT32), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(KEYINPUT32), .A3(new_n470), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n475));
  INV_X1    g289(.A(G119), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(G128), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n415), .A2(KEYINPUT23), .A3(G119), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n478), .C1(G119), .C2(new_n415), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G110), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT24), .B(G110), .Z(new_n481));
  XNOR2_X1  g295(.A(G119), .B(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n305), .B2(new_n312), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n479), .A2(G110), .B1(new_n482), .B2(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n293), .A2(new_n189), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n312), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT73), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT22), .B(G137), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(KEYINPUT74), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n485), .B2(new_n489), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n498), .B2(KEYINPUT75), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n381), .B1(G234), .B2(new_n281), .ZN(new_n503));
  INV_X1    g317(.A(new_n501), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n495), .A2(new_n497), .A3(new_n504), .A4(new_n499), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n497), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n503), .A2(G902), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT76), .Z(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G221), .B1(new_n380), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n190), .A2(new_n192), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n199), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n190), .A2(new_n192), .A3(new_n188), .A4(G128), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n252), .A2(new_n254), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n245), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n255), .B2(new_n422), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n411), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n252), .A2(new_n254), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n422), .B1(new_n245), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n518), .B1(new_n207), .B2(new_n416), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n253), .A2(KEYINPUT80), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n251), .B(new_n238), .C1(new_n231), .C2(new_n239), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n244), .B2(new_n242), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT12), .B(new_n411), .C1(new_n526), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n210), .A2(G227), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT77), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G140), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n236), .A2(new_n208), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n200), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n247), .A2(new_n539), .B1(new_n255), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n411), .B(KEYINPUT82), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n520), .B2(new_n540), .ZN(new_n545));
  AOI211_X1 g359(.A(KEYINPUT81), .B(KEYINPUT10), .C1(new_n245), .C2(new_n519), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n533), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n547), .ZN(new_n549));
  INV_X1    g363(.A(new_n411), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT83), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n542), .B(KEYINPUT83), .C1(new_n545), .C2(new_n546), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n548), .B1(new_n555), .B2(new_n538), .ZN(new_n556));
  OAI21_X1  g370(.A(G469), .B1(new_n556), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(G469), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT12), .B1(new_n521), .B2(new_n411), .ZN(new_n559));
  INV_X1    g373(.A(new_n532), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n547), .B(new_n537), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT84), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n533), .A2(KEYINPUT84), .A3(new_n537), .A4(new_n547), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n551), .A2(new_n552), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n411), .A3(new_n554), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n537), .B1(new_n567), .B2(new_n547), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n558), .B(new_n281), .C1(new_n565), .C2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n515), .B1(new_n557), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n397), .A2(new_n474), .A3(new_n513), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  INV_X1    g386(.A(G472), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n469), .B2(new_n281), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n470), .B2(new_n469), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n575), .A2(new_n570), .A3(new_n513), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT33), .B1(new_n384), .B2(new_n385), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n390), .A2(new_n578), .A3(new_n383), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n579), .A3(G478), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n391), .A2(new_n345), .A3(new_n281), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n345), .A2(new_n281), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n336), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n344), .B(new_n187), .C1(new_n278), .C2(new_n279), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  OR3_X1    g407(.A1(new_n332), .A2(new_n334), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n334), .A2(new_n593), .B1(G475), .B2(new_n320), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n587), .A2(new_n395), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n576), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  OR2_X1    g414(.A1(new_n496), .A2(KEYINPUT36), .ZN(new_n601));
  INV_X1    g415(.A(new_n490), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n510), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n506), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n187), .B(new_n606), .C1(new_n278), .C2(new_n279), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n396), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n575), .A3(new_n570), .A4(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT37), .B(G110), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n341), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n340), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n596), .A2(new_n395), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(new_n474), .A3(new_n570), .A4(new_n608), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  INV_X1    g433(.A(new_n473), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n471), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n281), .B1(new_n457), .B2(new_n441), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n442), .B1(new_n427), .B2(new_n434), .ZN(new_n623));
  OAI21_X1  g437(.A(G472), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT96), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n268), .A2(new_n276), .ZN(new_n628));
  INV_X1    g442(.A(new_n277), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n268), .A2(new_n276), .A3(new_n277), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n187), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n335), .A2(new_n394), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n606), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n615), .B(KEYINPUT39), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n570), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n627), .A2(new_n637), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT97), .B(G143), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G45));
  NAND2_X1  g458(.A1(new_n585), .A2(new_n615), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n474), .A3(new_n570), .A4(new_n608), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G146), .ZN(G48));
  NAND2_X1  g462(.A1(new_n474), .A2(new_n513), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n565), .A2(new_n568), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n281), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n652), .A3(G469), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n650), .B(new_n281), .C1(KEYINPUT98), .C2(new_n558), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n649), .A2(new_n655), .A3(new_n515), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n588), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G15));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n597), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  AOI21_X1  g475(.A(new_n635), .B1(new_n630), .B2(new_n631), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n653), .A2(new_n514), .A3(new_n662), .A4(new_n654), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n474), .A3(new_n609), .A4(new_n606), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  OAI211_X1 g480(.A(KEYINPUT99), .B(new_n468), .C1(new_n458), .C2(new_n441), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n466), .ZN(new_n668));
  INV_X1    g482(.A(new_n456), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n454), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n444), .B1(new_n670), .B2(new_n434), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n442), .B1(new_n671), .B2(new_n452), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT99), .B1(new_n672), .B2(new_n468), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n470), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n574), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(KEYINPUT100), .B(new_n470), .C1(new_n668), .C2(new_n673), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n655), .A2(new_n515), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n587), .A2(new_n636), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n513), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n363), .ZN(G24));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n606), .A3(new_n646), .A4(new_n677), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n663), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n201), .ZN(G27));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n630), .A2(new_n187), .A3(new_n631), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(G469), .A2(G902), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT101), .Z(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n556), .B2(G469), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n515), .B1(new_n691), .B2(new_n569), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g508(.A(KEYINPUT102), .B(new_n515), .C1(new_n691), .C2(new_n569), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n691), .A2(new_n569), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n514), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n692), .A2(new_n693), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(KEYINPUT103), .A3(new_n700), .A4(new_n688), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n649), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(KEYINPUT104), .B(KEYINPUT42), .C1(new_n702), .C2(new_n646), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n696), .A2(new_n701), .ZN(new_n705));
  INV_X1    g519(.A(new_n649), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n646), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n696), .B2(new_n701), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n620), .B2(new_n471), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n471), .A2(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .B1(G472), .B2(new_n461), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n717), .A3(new_n714), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n512), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n710), .B1(new_n712), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n712), .A2(new_n719), .A3(new_n710), .ZN(new_n721));
  OAI22_X1  g535(.A1(new_n703), .A2(new_n709), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT108), .B(G131), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G33));
  NAND2_X1  g538(.A1(new_n702), .A2(new_n617), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  AOI21_X1  g540(.A(new_n558), .B1(new_n556), .B2(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(KEYINPUT45), .B2(new_n556), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n690), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n569), .B1(new_n731), .B2(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n514), .B(new_n638), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n584), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n336), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT43), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT43), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n606), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n740), .A3(new_n575), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n740), .B1(new_n739), .B2(new_n575), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n688), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n734), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT110), .B(G137), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G39));
  OAI21_X1  g560(.A(new_n514), .B1(new_n732), .B2(new_n733), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT47), .B(new_n514), .C1(new_n732), .C2(new_n733), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n474), .A2(new_n645), .A3(new_n513), .A4(new_n687), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  NAND2_X1  g568(.A1(new_n626), .A2(new_n513), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n655), .A2(KEYINPUT49), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n655), .A2(KEYINPUT49), .ZN(new_n758));
  INV_X1    g572(.A(new_n634), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n759), .A2(new_n515), .A3(new_n635), .A4(new_n736), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n687), .A2(new_n340), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n626), .A2(new_n513), .A3(new_n679), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n735), .A2(new_n335), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n678), .A2(new_n606), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n679), .A2(new_n762), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n737), .A2(new_n738), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n340), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n513), .A3(new_n678), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n679), .A2(new_n635), .A3(new_n634), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT113), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n653), .A2(new_n515), .A3(new_n654), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n749), .A2(new_n750), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n772), .A2(new_n687), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n769), .A2(new_n719), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT48), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n338), .B1(new_n763), .B2(new_n586), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n772), .A2(new_n663), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n784), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n784), .B2(new_n788), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n782), .A2(KEYINPUT51), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n782), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n657), .A2(new_n660), .A3(new_n665), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(new_n681), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n649), .B(new_n645), .C1(new_n696), .C2(new_n701), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT104), .B1(new_n799), .B2(KEYINPUT42), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n707), .A2(new_n704), .A3(new_n708), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n712), .A2(new_n719), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT107), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n712), .A2(new_n719), .A3(new_n710), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n798), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n618), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n606), .A2(new_n676), .A3(new_n646), .A4(new_n677), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(new_n664), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n280), .A2(new_n606), .A3(new_n616), .A4(new_n636), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n625), .A3(new_n692), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n647), .A4(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n618), .B(new_n647), .C1(new_n683), .C2(new_n663), .ZN(new_n815));
  INV_X1    g629(.A(new_n813), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n335), .A2(new_n584), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n335), .B2(new_n394), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n587), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n513), .A3(new_n575), .A4(new_n570), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n606), .A2(new_n395), .A3(new_n615), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n687), .A2(new_n823), .A3(new_n596), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n474), .A3(new_n570), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n825), .A3(new_n571), .A4(new_n610), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n705), .B2(new_n809), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n725), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n807), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n798), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n810), .B2(new_n811), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n722), .A2(new_n829), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n722), .A2(new_n829), .A3(new_n831), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n832), .ZN(new_n838));
  INV_X1    g652(.A(new_n810), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n832), .B1(new_n839), .B2(KEYINPUT52), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n827), .A2(new_n725), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n827), .B2(new_n725), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n818), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n807), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n835), .A2(new_n836), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n836), .B1(new_n835), .B2(new_n848), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT116), .B(new_n796), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n337), .A2(new_n210), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n838), .A2(new_n846), .A3(new_n847), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n807), .A2(new_n829), .A3(new_n833), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n847), .B1(new_n838), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT112), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n835), .A2(new_n836), .A3(new_n848), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT116), .B1(new_n859), .B2(new_n796), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n761), .B1(new_n853), .B2(new_n860), .ZN(G75));
  NOR2_X1   g675(.A1(new_n210), .A2(G952), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT119), .Z(new_n863));
  AOI21_X1  g677(.A(new_n281), .B1(new_n838), .B2(new_n846), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n864), .B2(G210), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n272), .A2(new_n274), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n275), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n863), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n869), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G51));
  NAND2_X1  g688(.A1(new_n838), .A2(new_n846), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n848), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n690), .B(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n650), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n864), .A2(new_n730), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(G54));
  NAND3_X1  g698(.A1(new_n864), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  INV_X1    g699(.A(new_n330), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n862), .ZN(G60));
  AND2_X1   g703(.A1(new_n577), .A2(new_n579), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n583), .B(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n878), .A2(new_n879), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n863), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n849), .A2(new_n850), .A3(new_n892), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n890), .B2(new_n896), .ZN(G63));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n898));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n838), .B2(new_n846), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n603), .A3(new_n604), .ZN(new_n902));
  INV_X1    g716(.A(new_n863), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n875), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n507), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n907), .B(new_n863), .C1(new_n901), .C2(new_n508), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n898), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(KEYINPUT123), .A3(new_n507), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n901), .B2(new_n508), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n903), .A2(new_n898), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n912), .A2(new_n914), .A3(new_n902), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G66));
  AOI21_X1  g731(.A(new_n210), .B1(new_n343), .B2(G224), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n571), .A2(new_n831), .A3(new_n610), .A4(new_n822), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n210), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n866), .B1(G898), .B2(new_n210), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n921), .B(new_n922), .Z(G69));
  NOR4_X1   g737(.A1(new_n649), .A2(new_n639), .A3(new_n687), .A4(new_n820), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT124), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n744), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n642), .A2(new_n647), .A3(new_n810), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n753), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n210), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n426), .B(new_n325), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n210), .A2(G900), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n722), .A2(new_n725), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n719), .A2(new_n335), .A3(new_n394), .A4(new_n662), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n734), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n815), .B(new_n744), .C1(new_n751), .C2(new_n752), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n934), .B1(new_n942), .B2(new_n210), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n933), .B1(new_n943), .B2(new_n932), .ZN(new_n944));
  INV_X1    g758(.A(G227), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n945), .B2(new_n613), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n933), .C1(new_n943), .C2(new_n932), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n930), .B2(new_n920), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n862), .B1(new_n954), .B2(new_n623), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n435), .A2(new_n442), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n467), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n953), .B(new_n957), .C1(new_n830), .C2(new_n834), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n953), .B1(new_n942), .B2(new_n920), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n435), .A2(new_n441), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(G57));
endmodule


