

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759;

  INV_X2 U370 ( .A(G953), .ZN(n633) );
  XNOR2_X1 U371 ( .A(n515), .B(n514), .ZN(n555) );
  AND2_X1 U372 ( .A1(n435), .A2(n433), .ZN(n347) );
  OR2_X2 U373 ( .A1(n723), .A2(G902), .ZN(n515) );
  XNOR2_X2 U374 ( .A(n538), .B(n537), .ZN(n574) );
  XNOR2_X1 U375 ( .A(G116), .B(KEYINPUT3), .ZN(n457) );
  AND2_X1 U376 ( .A1(n402), .A2(n400), .ZN(n586) );
  AND2_X1 U377 ( .A1(n404), .A2(n350), .ZN(n402) );
  AND2_X1 U378 ( .A1(n436), .A2(n435), .ZN(n576) );
  AND2_X1 U379 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X1 U380 ( .A(n406), .B(KEYINPUT68), .ZN(n671) );
  XNOR2_X1 U381 ( .A(n382), .B(n457), .ZN(n519) );
  XNOR2_X1 U382 ( .A(n531), .B(n442), .ZN(n477) );
  XNOR2_X1 U383 ( .A(n741), .B(G101), .ZN(n525) );
  NAND2_X1 U384 ( .A1(n456), .A2(n455), .ZN(n382) );
  XNOR2_X1 U385 ( .A(n379), .B(G146), .ZN(n531) );
  XNOR2_X1 U386 ( .A(n498), .B(n451), .ZN(n741) );
  INV_X1 U387 ( .A(G113), .ZN(n454) );
  XOR2_X1 U388 ( .A(G107), .B(G110), .Z(n517) );
  XOR2_X1 U389 ( .A(G143), .B(G128), .Z(n498) );
  NOR2_X1 U390 ( .A1(n752), .A2(n759), .ZN(n559) );
  XNOR2_X1 U391 ( .A(n466), .B(G472), .ZN(n384) );
  NOR2_X1 U392 ( .A1(n640), .A2(G902), .ZN(n465) );
  NAND2_X1 U393 ( .A1(n386), .A2(n385), .ZN(n622) );
  XNOR2_X1 U394 ( .A(n609), .B(KEYINPUT6), .ZN(n619) );
  XNOR2_X1 U395 ( .A(n381), .B(n380), .ZN(n494) );
  XNOR2_X1 U396 ( .A(n445), .B(n450), .ZN(n381) );
  INV_X1 U397 ( .A(n739), .ZN(n380) );
  NAND2_X1 U398 ( .A1(n586), .A2(n662), .ZN(n703) );
  NAND2_X1 U399 ( .A1(n627), .A2(n626), .ZN(n395) );
  XNOR2_X1 U400 ( .A(n375), .B(n546), .ZN(n585) );
  XNOR2_X1 U401 ( .A(n505), .B(G478), .ZN(n562) );
  XOR2_X1 U402 ( .A(KEYINPUT91), .B(KEYINPUT94), .Z(n490) );
  XNOR2_X1 U403 ( .A(n469), .B(n468), .ZN(n491) );
  XNOR2_X1 U404 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n468) );
  INV_X1 U405 ( .A(G125), .ZN(n379) );
  INV_X1 U406 ( .A(n755), .ZN(n419) );
  NOR2_X1 U407 ( .A1(n425), .A2(n606), .ZN(n424) );
  OR2_X1 U408 ( .A1(n429), .A2(n754), .ZN(n426) );
  INV_X1 U409 ( .A(KEYINPUT77), .ZN(n575) );
  NOR2_X1 U410 ( .A1(n753), .A2(KEYINPUT44), .ZN(n626) );
  INV_X1 U411 ( .A(KEYINPUT22), .ZN(n596) );
  NOR2_X1 U412 ( .A1(n622), .A2(n595), .ZN(n597) );
  OR2_X1 U413 ( .A1(n684), .A2(n666), .ZN(n595) );
  XNOR2_X1 U414 ( .A(n464), .B(n463), .ZN(n640) );
  XOR2_X1 U415 ( .A(n504), .B(n503), .Z(n636) );
  XNOR2_X1 U416 ( .A(n525), .B(n452), .ZN(n508) );
  XNOR2_X1 U417 ( .A(n740), .B(G146), .ZN(n452) );
  NOR2_X1 U418 ( .A1(n568), .A2(n567), .ZN(n570) );
  AND2_X1 U419 ( .A1(n619), .A2(n618), .ZN(n621) );
  BUF_X1 U420 ( .A(n574), .Z(n568) );
  XNOR2_X1 U421 ( .A(n495), .B(n440), .ZN(n578) );
  BUF_X1 U422 ( .A(n622), .Z(n383) );
  XNOR2_X1 U423 ( .A(n488), .B(n487), .ZN(n637) );
  XNOR2_X1 U424 ( .A(n482), .B(n481), .ZN(n488) );
  INV_X1 U425 ( .A(n636), .ZN(n368) );
  NAND2_X1 U426 ( .A1(n371), .A2(n631), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n374), .A2(n373), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n508), .B(n411), .ZN(n723) );
  XNOR2_X1 U429 ( .A(n511), .B(n412), .ZN(n411) );
  XNOR2_X1 U430 ( .A(n512), .B(n509), .ZN(n412) );
  XNOR2_X1 U431 ( .A(n517), .B(n510), .ZN(n511) );
  OR2_X1 U432 ( .A1(n585), .A2(n660), .ZN(n662) );
  NOR2_X1 U433 ( .A1(n585), .A2(n657), .ZN(n548) );
  NOR2_X1 U434 ( .A1(n655), .A2(n580), .ZN(n581) );
  NAND2_X1 U435 ( .A1(n593), .A2(KEYINPUT0), .ZN(n433) );
  INV_X1 U436 ( .A(G119), .ZN(n453) );
  OR2_X1 U437 ( .A1(G902), .A2(G237), .ZN(n536) );
  XNOR2_X1 U438 ( .A(n399), .B(n492), .ZN(n418) );
  NAND2_X1 U439 ( .A1(n491), .A2(G217), .ZN(n399) );
  NAND2_X1 U440 ( .A1(n418), .A2(G902), .ZN(n416) );
  NAND2_X1 U441 ( .A1(n433), .A2(n594), .ZN(n430) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n446) );
  XNOR2_X1 U443 ( .A(n458), .B(n393), .ZN(n462) );
  XNOR2_X1 U444 ( .A(n459), .B(G131), .ZN(n393) );
  XOR2_X1 U445 ( .A(KEYINPUT9), .B(G116), .Z(n497) );
  XNOR2_X1 U446 ( .A(G122), .B(G107), .ZN(n496) );
  XNOR2_X1 U447 ( .A(n390), .B(n498), .ZN(n500) );
  XNOR2_X1 U448 ( .A(n499), .B(n391), .ZN(n390) );
  INV_X1 U449 ( .A(KEYINPUT7), .ZN(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT101), .B(G134), .ZN(n499) );
  XOR2_X1 U451 ( .A(G134), .B(G137), .Z(n740) );
  XNOR2_X1 U452 ( .A(KEYINPUT87), .B(KEYINPUT79), .ZN(n528) );
  NAND2_X1 U453 ( .A1(n401), .A2(KEYINPUT48), .ZN(n400) );
  NAND2_X1 U454 ( .A1(n432), .A2(n351), .ZN(n435) );
  NAND2_X1 U455 ( .A1(n605), .A2(n407), .ZN(n406) );
  INV_X1 U456 ( .A(n666), .ZN(n407) );
  XNOR2_X1 U457 ( .A(G128), .B(G137), .ZN(n484) );
  XNOR2_X1 U458 ( .A(n423), .B(n422), .ZN(n480) );
  XNOR2_X1 U459 ( .A(KEYINPUT23), .B(G140), .ZN(n423) );
  XNOR2_X1 U460 ( .A(G110), .B(G119), .ZN(n422) );
  XNOR2_X1 U461 ( .A(G902), .B(KEYINPUT15), .ZN(n630) );
  XNOR2_X1 U462 ( .A(G140), .B(G131), .ZN(n512) );
  INV_X1 U463 ( .A(G104), .ZN(n509) );
  NAND2_X1 U464 ( .A1(G237), .A2(G234), .ZN(n473) );
  NOR2_X1 U465 ( .A1(n609), .A2(n573), .ZN(n541) );
  NOR2_X1 U466 ( .A1(n557), .A2(n556), .ZN(n577) );
  XNOR2_X1 U467 ( .A(n398), .B(KEYINPUT67), .ZN(n429) );
  XNOR2_X1 U468 ( .A(n572), .B(KEYINPUT110), .ZN(n756) );
  XNOR2_X1 U469 ( .A(n408), .B(KEYINPUT35), .ZN(n753) );
  XNOR2_X1 U470 ( .A(n428), .B(KEYINPUT32), .ZN(n427) );
  INV_X1 U471 ( .A(KEYINPUT66), .ZN(n428) );
  AND2_X1 U472 ( .A1(n429), .A2(n598), .ZN(n650) );
  INV_X1 U473 ( .A(n562), .ZN(n579) );
  INV_X1 U474 ( .A(n578), .ZN(n389) );
  NOR2_X1 U475 ( .A1(n614), .A2(n667), .ZN(n615) );
  XNOR2_X1 U476 ( .A(n358), .B(n356), .ZN(G57) );
  XNOR2_X1 U477 ( .A(n377), .B(n376), .ZN(n392) );
  INV_X1 U478 ( .A(n637), .ZN(n376) );
  XNOR2_X1 U479 ( .A(n362), .B(n361), .ZN(G63) );
  INV_X1 U480 ( .A(KEYINPUT122), .ZN(n361) );
  XNOR2_X1 U481 ( .A(n360), .B(n359), .ZN(G60) );
  INV_X1 U482 ( .A(KEYINPUT60), .ZN(n359) );
  XNOR2_X1 U483 ( .A(n721), .B(n387), .ZN(n724) );
  XNOR2_X1 U484 ( .A(n723), .B(n722), .ZN(n387) );
  AND2_X1 U485 ( .A1(n662), .A2(KEYINPUT2), .ZN(n348) );
  XOR2_X1 U486 ( .A(n575), .B(KEYINPUT19), .Z(n349) );
  XNOR2_X1 U487 ( .A(n465), .B(n384), .ZN(n674) );
  INV_X1 U488 ( .A(n674), .ZN(n609) );
  AND2_X1 U489 ( .A1(n403), .A2(n419), .ZN(n350) );
  OR2_X1 U490 ( .A1(n413), .A2(n415), .ZN(n605) );
  INV_X1 U491 ( .A(n593), .ZN(n434) );
  NOR2_X1 U492 ( .A1(n573), .A2(n349), .ZN(n351) );
  INV_X1 U493 ( .A(n605), .ZN(n598) );
  AND2_X1 U494 ( .A1(n434), .A2(n594), .ZN(n352) );
  INV_X1 U495 ( .A(KEYINPUT0), .ZN(n594) );
  XOR2_X1 U496 ( .A(KEYINPUT82), .B(KEYINPUT45), .Z(n353) );
  XNOR2_X1 U497 ( .A(n494), .B(KEYINPUT59), .ZN(n354) );
  INV_X1 U498 ( .A(KEYINPUT2), .ZN(n629) );
  XOR2_X1 U499 ( .A(n640), .B(n639), .Z(n355) );
  XNOR2_X1 U500 ( .A(KEYINPUT86), .B(n634), .ZN(n725) );
  INV_X1 U501 ( .A(n725), .ZN(n366) );
  XOR2_X1 U502 ( .A(KEYINPUT85), .B(KEYINPUT63), .Z(n356) );
  XNOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n357) );
  NAND2_X1 U504 ( .A1(n364), .A2(n366), .ZN(n358) );
  NAND2_X1 U505 ( .A1(n365), .A2(n366), .ZN(n360) );
  NAND2_X1 U506 ( .A1(n367), .A2(n366), .ZN(n362) );
  XNOR2_X1 U507 ( .A(n363), .B(n357), .ZN(G51) );
  NAND2_X1 U508 ( .A1(n719), .A2(n366), .ZN(n363) );
  XNOR2_X1 U509 ( .A(n641), .B(n355), .ZN(n364) );
  XNOR2_X1 U510 ( .A(n632), .B(n354), .ZN(n365) );
  XNOR2_X1 U511 ( .A(n635), .B(n368), .ZN(n367) );
  OR2_X2 U512 ( .A1(n369), .A2(n734), .ZN(n374) );
  XNOR2_X2 U513 ( .A(n394), .B(n353), .ZN(n734) );
  NAND2_X1 U514 ( .A1(n586), .A2(n348), .ZN(n369) );
  NOR2_X1 U515 ( .A1(n703), .A2(n734), .ZN(n705) );
  NOR2_X4 U516 ( .A1(n372), .A2(n370), .ZN(n720) );
  NAND2_X1 U517 ( .A1(n734), .A2(n629), .ZN(n371) );
  NAND2_X1 U518 ( .A1(n703), .A2(n629), .ZN(n373) );
  NAND2_X1 U519 ( .A1(n561), .A2(n545), .ZN(n375) );
  NOR2_X1 U520 ( .A1(n607), .A2(n543), .ZN(n544) );
  XNOR2_X1 U521 ( .A(n542), .B(KEYINPUT95), .ZN(n607) );
  NAND2_X1 U522 ( .A1(n720), .A2(G217), .ZN(n377) );
  BUF_X1 U523 ( .A(n726), .Z(n378) );
  NAND2_X1 U524 ( .A1(n720), .A2(G478), .ZN(n635) );
  XNOR2_X1 U525 ( .A(n522), .B(n521), .ZN(n726) );
  NAND2_X1 U526 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U527 ( .A1(n642), .A2(n616), .ZN(n617) );
  NAND2_X1 U528 ( .A1(n615), .A2(n670), .ZN(n642) );
  NAND2_X1 U529 ( .A1(n576), .A2(n352), .ZN(n385) );
  NAND2_X1 U530 ( .A1(n431), .A2(n430), .ZN(n386) );
  XNOR2_X1 U531 ( .A(n397), .B(KEYINPUT65), .ZN(n396) );
  NOR2_X1 U532 ( .A1(n396), .A2(n628), .ZN(n388) );
  NOR2_X1 U533 ( .A1(n663), .A2(n383), .ZN(n410) );
  NAND2_X1 U534 ( .A1(n388), .A2(n395), .ZN(n394) );
  NOR2_X1 U535 ( .A1(n754), .A2(n598), .ZN(n425) );
  NAND2_X1 U536 ( .A1(n562), .A2(n389), .ZN(n657) );
  NAND2_X1 U537 ( .A1(n392), .A2(n366), .ZN(n638) );
  NAND2_X1 U538 ( .A1(n426), .A2(n424), .ZN(n397) );
  NAND2_X1 U539 ( .A1(n604), .A2(n609), .ZN(n398) );
  INV_X1 U540 ( .A(n566), .ZN(n401) );
  OR2_X1 U541 ( .A1(n420), .A2(n584), .ZN(n403) );
  NAND2_X1 U542 ( .A1(n566), .A2(n405), .ZN(n404) );
  AND2_X1 U543 ( .A1(n420), .A2(n584), .ZN(n405) );
  NAND2_X1 U544 ( .A1(n409), .A2(n623), .ZN(n408) );
  XNOR2_X1 U545 ( .A(n410), .B(KEYINPUT34), .ZN(n409) );
  NOR2_X1 U546 ( .A1(n637), .A2(n414), .ZN(n413) );
  OR2_X1 U547 ( .A1(n418), .A2(G902), .ZN(n414) );
  NAND2_X1 U548 ( .A1(n637), .A2(n418), .ZN(n417) );
  NOR2_X1 U549 ( .A1(n583), .A2(n421), .ZN(n420) );
  INV_X1 U550 ( .A(n654), .ZN(n421) );
  XNOR2_X2 U551 ( .A(n600), .B(n427), .ZN(n754) );
  NOR2_X1 U552 ( .A1(n650), .A2(n754), .ZN(n627) );
  NAND2_X1 U553 ( .A1(n347), .A2(n436), .ZN(n431) );
  INV_X1 U554 ( .A(n574), .ZN(n432) );
  NAND2_X1 U555 ( .A1(n573), .A2(n349), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n574), .A2(n349), .ZN(n438) );
  XNOR2_X1 U557 ( .A(n597), .B(n596), .ZN(n601) );
  XOR2_X1 U558 ( .A(n448), .B(n447), .Z(n439) );
  XOR2_X1 U559 ( .A(KEYINPUT13), .B(G475), .Z(n440) );
  XNOR2_X1 U560 ( .A(n441), .B(KEYINPUT10), .ZN(n442) );
  NAND2_X1 U561 ( .A1(n578), .A2(n562), .ZN(n684) );
  XNOR2_X1 U562 ( .A(n480), .B(KEYINPUT78), .ZN(n481) );
  XNOR2_X1 U563 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U564 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U565 ( .A1(n555), .A2(n671), .ZN(n542) );
  XNOR2_X1 U566 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U567 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n546) );
  XNOR2_X1 U568 ( .A(n718), .B(n717), .ZN(n719) );
  INV_X1 U569 ( .A(n512), .ZN(n443) );
  INV_X1 U570 ( .A(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U571 ( .A(n443), .B(n477), .ZN(n739) );
  XOR2_X1 U572 ( .A(G122), .B(G104), .Z(n520) );
  XNOR2_X1 U573 ( .A(G143), .B(n520), .ZN(n444) );
  XNOR2_X1 U574 ( .A(n444), .B(G113), .ZN(n445) );
  XOR2_X1 U575 ( .A(KEYINPUT75), .B(n446), .Z(n460) );
  NAND2_X1 U576 ( .A1(n460), .A2(G214), .ZN(n449) );
  XOR2_X1 U577 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n448) );
  XNOR2_X1 U578 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n447) );
  XNOR2_X1 U579 ( .A(n449), .B(n439), .ZN(n450) );
  XNOR2_X1 U580 ( .A(KEYINPUT74), .B(KEYINPUT97), .ZN(n466) );
  XOR2_X1 U581 ( .A(KEYINPUT64), .B(KEYINPUT4), .Z(n451) );
  INV_X1 U582 ( .A(n508), .ZN(n464) );
  XOR2_X1 U583 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n459) );
  NAND2_X1 U584 ( .A1(G113), .A2(n453), .ZN(n456) );
  NAND2_X1 U585 ( .A1(n454), .A2(G119), .ZN(n455) );
  BUF_X1 U586 ( .A(n519), .Z(n458) );
  NAND2_X1 U587 ( .A1(G210), .A2(n460), .ZN(n461) );
  NAND2_X1 U588 ( .A1(n536), .A2(G214), .ZN(n467) );
  XOR2_X1 U589 ( .A(KEYINPUT88), .B(n467), .Z(n573) );
  INV_X1 U590 ( .A(n573), .ZN(n686) );
  NAND2_X1 U591 ( .A1(n630), .A2(G234), .ZN(n469) );
  NAND2_X1 U592 ( .A1(n491), .A2(G221), .ZN(n470) );
  XNOR2_X1 U593 ( .A(KEYINPUT21), .B(n470), .ZN(n666) );
  NOR2_X1 U594 ( .A1(G900), .A2(n633), .ZN(n471) );
  NAND2_X1 U595 ( .A1(n471), .A2(G902), .ZN(n472) );
  NAND2_X1 U596 ( .A1(G952), .A2(n633), .ZN(n590) );
  NAND2_X1 U597 ( .A1(n472), .A2(n590), .ZN(n474) );
  XNOR2_X1 U598 ( .A(n473), .B(KEYINPUT14), .ZN(n665) );
  NAND2_X1 U599 ( .A1(n474), .A2(n665), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n666), .A2(n543), .ZN(n493) );
  INV_X1 U601 ( .A(n477), .ZN(n475) );
  NAND2_X1 U602 ( .A1(n475), .A2(KEYINPUT24), .ZN(n479) );
  INV_X1 U603 ( .A(KEYINPUT24), .ZN(n476) );
  NAND2_X1 U604 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U605 ( .A1(n479), .A2(n478), .ZN(n482) );
  NAND2_X1 U606 ( .A1(G234), .A2(n633), .ZN(n483) );
  XOR2_X1 U607 ( .A(KEYINPUT8), .B(n483), .Z(n502) );
  NAND2_X1 U608 ( .A1(G221), .A2(n502), .ZN(n486) );
  XNOR2_X1 U609 ( .A(n484), .B(KEYINPUT80), .ZN(n485) );
  XNOR2_X1 U610 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n489) );
  XNOR2_X1 U611 ( .A(n490), .B(n489), .ZN(n492) );
  NAND2_X1 U612 ( .A1(n493), .A2(n598), .ZN(n552) );
  NOR2_X1 U613 ( .A1(G902), .A2(n494), .ZN(n495) );
  XNOR2_X1 U614 ( .A(n497), .B(n496), .ZN(n501) );
  XOR2_X1 U615 ( .A(n501), .B(n500), .Z(n504) );
  NAND2_X1 U616 ( .A1(G217), .A2(n502), .ZN(n503) );
  NOR2_X1 U617 ( .A1(G902), .A2(n636), .ZN(n505) );
  NOR2_X1 U618 ( .A1(n552), .A2(n657), .ZN(n506) );
  AND2_X1 U619 ( .A1(n686), .A2(n506), .ZN(n507) );
  NAND2_X1 U620 ( .A1(n619), .A2(n507), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G227), .A2(n633), .ZN(n510) );
  XNOR2_X1 U622 ( .A(G469), .B(KEYINPUT70), .ZN(n513) );
  XNOR2_X1 U623 ( .A(n513), .B(KEYINPUT71), .ZN(n514) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT1), .ZN(n670) );
  INV_X1 U625 ( .A(n670), .ZN(n602) );
  OR2_X1 U626 ( .A1(n567), .A2(n602), .ZN(n516) );
  XNOR2_X1 U627 ( .A(n516), .B(KEYINPUT43), .ZN(n539) );
  INV_X1 U628 ( .A(n517), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n519), .B(n518), .ZN(n522) );
  XNOR2_X1 U630 ( .A(KEYINPUT16), .B(n520), .ZN(n521) );
  INV_X1 U631 ( .A(n726), .ZN(n524) );
  INV_X1 U632 ( .A(n525), .ZN(n523) );
  NAND2_X1 U633 ( .A1(n524), .A2(n523), .ZN(n527) );
  NAND2_X1 U634 ( .A1(n726), .A2(n525), .ZN(n526) );
  NAND2_X1 U635 ( .A1(n527), .A2(n526), .ZN(n535) );
  XOR2_X1 U636 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n529) );
  XNOR2_X1 U637 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U638 ( .A(n531), .B(n530), .Z(n533) );
  NAND2_X1 U639 ( .A1(G224), .A2(n633), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U641 ( .A(n535), .B(n534), .ZN(n714) );
  NAND2_X1 U642 ( .A1(n714), .A2(n630), .ZN(n538) );
  NAND2_X1 U643 ( .A1(G210), .A2(n536), .ZN(n537) );
  NAND2_X1 U644 ( .A1(n539), .A2(n568), .ZN(n540) );
  XNOR2_X1 U645 ( .A(KEYINPUT105), .B(n540), .ZN(n755) );
  INV_X1 U646 ( .A(KEYINPUT48), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT30), .B(n541), .ZN(n560) );
  XNOR2_X1 U648 ( .A(KEYINPUT38), .B(n568), .ZN(n682) );
  AND2_X1 U649 ( .A1(n560), .A2(n682), .ZN(n545) );
  XNOR2_X1 U650 ( .A(n544), .B(KEYINPUT76), .ZN(n561) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n547) );
  XNOR2_X1 U652 ( .A(n548), .B(n547), .ZN(n752) );
  INV_X1 U653 ( .A(n684), .ZN(n549) );
  NAND2_X1 U654 ( .A1(n682), .A2(n549), .ZN(n689) );
  NOR2_X1 U655 ( .A1(n573), .A2(n689), .ZN(n551) );
  XNOR2_X1 U656 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n550) );
  XNOR2_X1 U657 ( .A(n551), .B(n550), .ZN(n681) );
  XOR2_X1 U658 ( .A(KEYINPUT107), .B(KEYINPUT28), .Z(n554) );
  OR2_X1 U659 ( .A1(n552), .A2(n609), .ZN(n553) );
  XNOR2_X1 U660 ( .A(n554), .B(n553), .ZN(n557) );
  XNOR2_X1 U661 ( .A(KEYINPUT106), .B(n555), .ZN(n556) );
  NAND2_X1 U662 ( .A1(n681), .A2(n577), .ZN(n558) );
  XOR2_X1 U663 ( .A(KEYINPUT42), .B(n558), .Z(n759) );
  XNOR2_X1 U664 ( .A(n559), .B(KEYINPUT46), .ZN(n566) );
  AND2_X1 U665 ( .A1(n561), .A2(n560), .ZN(n565) );
  NOR2_X1 U666 ( .A1(n578), .A2(n562), .ZN(n623) );
  INV_X1 U667 ( .A(n623), .ZN(n563) );
  NOR2_X1 U668 ( .A1(n568), .A2(n563), .ZN(n564) );
  NAND2_X1 U669 ( .A1(n565), .A2(n564), .ZN(n654) );
  XNOR2_X1 U670 ( .A(KEYINPUT36), .B(KEYINPUT84), .ZN(n569) );
  XNOR2_X1 U671 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U672 ( .A1(n571), .A2(n602), .ZN(n572) );
  NAND2_X1 U673 ( .A1(n577), .A2(n576), .ZN(n655) );
  NAND2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n660) );
  NAND2_X1 U675 ( .A1(n657), .A2(n660), .ZN(n683) );
  INV_X1 U676 ( .A(n683), .ZN(n580) );
  XNOR2_X1 U677 ( .A(n581), .B(KEYINPUT47), .ZN(n582) );
  NAND2_X1 U678 ( .A1(n756), .A2(n582), .ZN(n583) );
  XNOR2_X1 U679 ( .A(G898), .B(KEYINPUT89), .ZN(n732) );
  NAND2_X1 U680 ( .A1(G953), .A2(n732), .ZN(n729) );
  NAND2_X1 U681 ( .A1(G902), .A2(n665), .ZN(n587) );
  NOR2_X1 U682 ( .A1(n729), .A2(n587), .ZN(n588) );
  XNOR2_X1 U683 ( .A(n588), .B(KEYINPUT90), .ZN(n592) );
  INV_X1 U684 ( .A(n665), .ZN(n589) );
  NOR2_X1 U685 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U687 ( .A1(n601), .A2(n619), .ZN(n613) );
  XNOR2_X1 U688 ( .A(KEYINPUT102), .B(n598), .ZN(n667) );
  AND2_X1 U689 ( .A1(n602), .A2(n667), .ZN(n599) );
  NAND2_X1 U690 ( .A1(n613), .A2(n599), .ZN(n600) );
  NOR2_X1 U691 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U692 ( .A(n603), .B(KEYINPUT104), .ZN(n604) );
  INV_X1 U693 ( .A(KEYINPUT44), .ZN(n606) );
  NOR2_X1 U694 ( .A1(n383), .A2(n607), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n644) );
  NOR2_X1 U696 ( .A1(n671), .A2(n670), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n674), .A2(n618), .ZN(n610) );
  XNOR2_X1 U698 ( .A(n610), .B(KEYINPUT98), .ZN(n678) );
  NOR2_X1 U699 ( .A1(n678), .A2(n383), .ZN(n611) );
  XNOR2_X1 U700 ( .A(n611), .B(KEYINPUT31), .ZN(n659) );
  NAND2_X1 U701 ( .A1(n644), .A2(n659), .ZN(n612) );
  NAND2_X1 U702 ( .A1(n612), .A2(n683), .ZN(n616) );
  XNOR2_X1 U703 ( .A(KEYINPUT83), .B(n613), .ZN(n614) );
  XNOR2_X1 U704 ( .A(n617), .B(KEYINPUT103), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n620) );
  XNOR2_X1 U706 ( .A(n621), .B(n620), .ZN(n663) );
  NAND2_X1 U707 ( .A1(KEYINPUT44), .A2(n753), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n628) );
  INV_X1 U709 ( .A(n630), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n720), .A2(G475), .ZN(n632) );
  NOR2_X1 U711 ( .A1(G952), .A2(n633), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n638), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U713 ( .A1(n720), .A2(G472), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT62), .B(KEYINPUT111), .Z(n639) );
  XNOR2_X1 U715 ( .A(G101), .B(n642), .ZN(G3) );
  NOR2_X1 U716 ( .A1(n657), .A2(n644), .ZN(n643) );
  XOR2_X1 U717 ( .A(G104), .B(n643), .Z(G6) );
  NOR2_X1 U718 ( .A1(n660), .A2(n644), .ZN(n649) );
  XOR2_X1 U719 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n646) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT26), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT27), .B(n647), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(G9) );
  XOR2_X1 U724 ( .A(G110), .B(n650), .Z(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT114), .B(n651), .ZN(G12) );
  NOR2_X1 U726 ( .A1(n660), .A2(n655), .ZN(n653) );
  XNOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(G30) );
  XNOR2_X1 U729 ( .A(G143), .B(n654), .ZN(G45) );
  NOR2_X1 U730 ( .A1(n657), .A2(n655), .ZN(n656) );
  XOR2_X1 U731 ( .A(G146), .B(n656), .Z(G48) );
  NOR2_X1 U732 ( .A1(n657), .A2(n659), .ZN(n658) );
  XOR2_X1 U733 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U735 ( .A(G116), .B(n661), .Z(G18) );
  XNOR2_X1 U736 ( .A(G134), .B(n662), .ZN(G36) );
  INV_X1 U737 ( .A(n663), .ZN(n691) );
  AND2_X1 U738 ( .A1(n691), .A2(n681), .ZN(n664) );
  NOR2_X1 U739 ( .A1(G953), .A2(n664), .ZN(n702) );
  NAND2_X1 U740 ( .A1(G952), .A2(n665), .ZN(n699) );
  XNOR2_X1 U741 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n697) );
  XOR2_X1 U742 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n669) );
  NAND2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n669), .B(n668), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U746 ( .A(KEYINPUT50), .B(n672), .Z(n673) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NAND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U756 ( .A(KEYINPUT117), .B(n690), .Z(n692) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n695), .B(KEYINPUT52), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U762 ( .A(KEYINPUT120), .B(n700), .Z(n701) );
  NAND2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n712) );
  INV_X1 U764 ( .A(n703), .ZN(n744) );
  NOR2_X1 U765 ( .A1(KEYINPUT2), .A2(n744), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n704), .B(KEYINPUT81), .ZN(n707) );
  NAND2_X1 U767 ( .A1(KEYINPUT2), .A2(n705), .ZN(n706) );
  NAND2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n710) );
  INV_X1 U769 ( .A(n734), .ZN(n708) );
  NOR2_X1 U770 ( .A1(KEYINPUT2), .A2(n708), .ZN(n709) );
  NOR2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U773 ( .A(KEYINPUT53), .B(n713), .ZN(G75) );
  NAND2_X1 U774 ( .A1(n720), .A2(G210), .ZN(n718) );
  BUF_X1 U775 ( .A(n714), .Z(n716) );
  XOR2_X1 U776 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n715) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n722) );
  NAND2_X1 U778 ( .A1(n720), .A2(G469), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n725), .A2(n724), .ZN(G54) );
  XNOR2_X1 U780 ( .A(G101), .B(n378), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n727), .B(KEYINPUT125), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n738) );
  XOR2_X1 U783 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n731) );
  NAND2_X1 U784 ( .A1(G224), .A2(G953), .ZN(n730) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U787 ( .A1(G953), .A2(n734), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT126), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n747), .B(n744), .ZN(n745) );
  NOR2_X1 U794 ( .A1(G953), .A2(n745), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n746), .B(KEYINPUT127), .ZN(n751) );
  XNOR2_X1 U796 ( .A(G227), .B(n747), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U800 ( .A(G131), .B(n752), .Z(G33) );
  XOR2_X1 U801 ( .A(G122), .B(n753), .Z(G24) );
  XOR2_X1 U802 ( .A(G119), .B(n754), .Z(G21) );
  XOR2_X1 U803 ( .A(G140), .B(n755), .Z(G42) );
  XNOR2_X1 U804 ( .A(n756), .B(KEYINPUT115), .ZN(n757) );
  XNOR2_X1 U805 ( .A(n757), .B(KEYINPUT37), .ZN(n758) );
  XNOR2_X1 U806 ( .A(G125), .B(n758), .ZN(G27) );
  XOR2_X1 U807 ( .A(n759), .B(G137), .Z(G39) );
endmodule

