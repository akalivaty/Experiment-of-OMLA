//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n191), .A3(G143), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n193), .B(G146), .C1(new_n203), .C2(KEYINPUT1), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n205), .C1(new_n195), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n202), .B1(G125), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G224), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(KEYINPUT5), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT74), .A2(G104), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT74), .A2(G104), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT74), .A2(G104), .ZN(new_n235));
  OAI21_X1  g049(.A(G107), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT75), .A2(G107), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT75), .A2(G107), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n232), .A2(new_n233), .A3(new_n236), .A4(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT75), .B(G107), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n231), .B1(new_n242), .B2(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n241), .B2(new_n244), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n219), .B(new_n225), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT80), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT76), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n219), .A4(new_n225), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n234), .A2(new_n235), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n229), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n240), .A2(new_n236), .ZN(new_n259));
  OAI21_X1  g073(.A(G101), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n261));
  INV_X1    g075(.A(G119), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G116), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n214), .B(new_n216), .C1(new_n222), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n219), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G101), .C1(new_n258), .C2(new_n259), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n249), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  XOR2_X1   g084(.A(G110), .B(G122), .Z(new_n271));
  NAND4_X1  g085(.A1(new_n269), .A2(KEYINPUT81), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n269), .A2(KEYINPUT81), .A3(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT6), .B1(new_n269), .B2(new_n271), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n212), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n211), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n212), .B(new_n279), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n271), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n220), .A3(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n219), .B(new_n285), .C1(new_n246), .C2(new_n247), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n253), .A2(KEYINPUT83), .A3(new_n219), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n225), .A2(new_n219), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n288), .A2(new_n289), .B1(new_n250), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT8), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n282), .B(new_n269), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n271), .B1(new_n291), .B2(KEYINPUT8), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n190), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n294), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n280), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(new_n276), .A3(new_n189), .A4(new_n275), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G475), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n304), .A2(KEYINPUT16), .A3(G140), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(KEYINPUT16), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n191), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G214), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n193), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(G143), .A3(G214), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT17), .ZN(new_n315));
  INV_X1    g129(.A(new_n313), .ZN(new_n316));
  AOI21_X1  g130(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n317));
  OAI21_X1  g131(.A(G131), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n312), .A2(new_n309), .A3(new_n313), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n308), .B(new_n315), .C1(KEYINPUT17), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(KEYINPUT18), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n316), .A2(new_n317), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n306), .A2(new_n191), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n191), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G113), .B(G122), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(new_n227), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT87), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n330), .B2(new_n333), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n303), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n306), .A2(KEYINPUT85), .A3(KEYINPUT19), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT19), .B1(new_n306), .B2(KEYINPUT85), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n191), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n318), .A2(new_n319), .B1(G146), .B2(new_n307), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n323), .A2(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n322), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n337), .B1(new_n344), .B2(new_n332), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n329), .ZN(new_n347));
  INV_X1    g161(.A(new_n332), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(KEYINPUT86), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n321), .A2(new_n332), .A3(new_n329), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n303), .A3(new_n276), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT20), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n351), .A2(new_n354), .A3(new_n303), .A4(new_n276), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n336), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G128), .B(G143), .ZN(new_n357));
  INV_X1    g171(.A(G134), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G116), .B(G122), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n242), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT14), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n221), .A2(KEYINPUT14), .A3(G122), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(G107), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n203), .A2(KEYINPUT13), .A3(G143), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n358), .B(new_n367), .C1(KEYINPUT13), .C2(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n357), .A2(new_n358), .ZN(new_n369));
  INV_X1    g183(.A(new_n361), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n242), .A2(new_n360), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n366), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT9), .B(G234), .Z(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(G217), .A3(new_n210), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT88), .Z(new_n376));
  OR2_X1    g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n376), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G478), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT15), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n379), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n210), .A2(G952), .ZN(new_n384));
  NAND2_X1  g198(.A1(G234), .A2(G237), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n386), .B(KEYINPUT89), .Z(new_n387));
  XOR2_X1   g201(.A(KEYINPUT21), .B(G898), .Z(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(G902), .A3(G953), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n356), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n300), .A2(new_n302), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n203), .A2(G119), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n393), .A2(KEYINPUT72), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n262), .A2(G128), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT72), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n308), .B1(G110), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n203), .A2(KEYINPUT69), .A3(G119), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT69), .B1(new_n203), .B2(G119), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT24), .B(G110), .Z(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n403), .B(KEYINPUT70), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT71), .A3(new_n407), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n400), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n307), .A2(G146), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(new_n407), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n399), .A2(G110), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n414), .B(new_n327), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT22), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(G137), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n413), .B2(new_n417), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT25), .A3(new_n276), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n413), .A2(new_n417), .ZN(new_n426));
  INV_X1    g240(.A(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n276), .A3(new_n421), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G217), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(G234), .B2(new_n276), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n424), .A2(new_n276), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n310), .A2(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n233), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(new_n233), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT26), .B(KEYINPUT27), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G101), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(G210), .A3(new_n310), .A4(new_n441), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT11), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n358), .B2(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n358), .A2(G137), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT11), .A3(G134), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G131), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n450), .A2(new_n453), .A3(new_n309), .A4(new_n451), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n201), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(KEYINPUT64), .A3(G134), .ZN(new_n459));
  INV_X1    g273(.A(new_n451), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT64), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n358), .B2(G137), .ZN(new_n462));
  OAI211_X1 g276(.A(G131), .B(new_n459), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n207), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n264), .A2(new_n219), .A3(KEYINPUT65), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT65), .B1(new_n264), .B2(new_n219), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n448), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n464), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n455), .A2(new_n456), .B1(new_n199), .B2(new_n200), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT30), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n458), .B2(new_n464), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n265), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n458), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT66), .A3(new_n448), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT31), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n471), .A2(new_n477), .A3(KEYINPUT31), .A4(new_n479), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n265), .B1(new_n472), .B2(new_n473), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n484), .A3(KEYINPUT67), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n465), .A2(new_n486), .A3(new_n265), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(KEYINPUT28), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n478), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n448), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n482), .A2(new_n483), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(G472), .A2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(KEYINPUT68), .B(KEYINPUT32), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n482), .A2(new_n483), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n492), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n494), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n493), .B2(new_n495), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n497), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n477), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(new_n489), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n492), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n492), .C2(new_n491), .ZN(new_n513));
  INV_X1    g327(.A(new_n490), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n465), .A2(new_n468), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n478), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n516), .B2(KEYINPUT28), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n492), .A2(new_n512), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G472), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n438), .B1(new_n507), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G221), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n374), .B2(new_n276), .ZN(new_n524));
  INV_X1    g338(.A(G469), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n246), .A2(new_n247), .A3(new_n207), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n250), .A2(new_n208), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n457), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(KEYINPUT78), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(KEYINPUT78), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n261), .A2(new_n201), .A3(new_n267), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n250), .B2(new_n208), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT10), .B(new_n207), .C1(new_n246), .C2(new_n247), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT77), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n253), .A2(new_n539), .A3(KEYINPUT10), .A4(new_n207), .ZN(new_n540));
  INV_X1    g354(.A(new_n457), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n527), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n253), .B2(new_n207), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT78), .A3(new_n529), .A4(new_n457), .ZN(new_n545));
  XOR2_X1   g359(.A(G110), .B(G140), .Z(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  INV_X1    g361(.A(G227), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G953), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n547), .B(new_n549), .Z(new_n550));
  NAND4_X1  g364(.A1(new_n532), .A2(new_n542), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n538), .A2(new_n536), .A3(new_n540), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n457), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n554), .B2(new_n542), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n525), .B(new_n276), .C1(new_n552), .C2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT79), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n542), .ZN(new_n559));
  INV_X1    g373(.A(new_n550), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n551), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(KEYINPUT79), .A3(new_n525), .A4(new_n276), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n554), .A2(new_n542), .A3(new_n550), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n532), .A2(new_n542), .A3(new_n545), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n276), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G469), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n524), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n392), .A2(new_n522), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n277), .B2(new_n295), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n298), .A2(KEYINPUT91), .A3(new_n276), .A4(new_n275), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n574), .A2(new_n188), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n573), .B(new_n187), .C1(new_n277), .C2(new_n295), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n301), .ZN(new_n578));
  INV_X1    g392(.A(new_n390), .ZN(new_n579));
  INV_X1    g393(.A(new_n378), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT33), .B1(new_n580), .B2(KEYINPUT92), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n377), .A2(new_n378), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n377), .A2(KEYINPUT92), .A3(KEYINPUT33), .A4(new_n378), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(new_n584), .A3(G478), .A4(new_n276), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT93), .B(G478), .Z(new_n586));
  OR2_X1    g400(.A1(new_n379), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n356), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n561), .B2(new_n551), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT79), .B1(new_n592), .B2(new_n525), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n556), .A2(new_n557), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n569), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n438), .A2(new_n524), .ZN(new_n596));
  OAI21_X1  g410(.A(G472), .B1(new_n493), .B2(G902), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n505), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n595), .A2(KEYINPUT90), .A3(new_n596), .A4(new_n598), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n591), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(new_n355), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n336), .B1(new_n606), .B2(KEYINPUT94), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n353), .A2(new_n608), .A3(new_n355), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n609), .A3(new_n382), .ZN(new_n610));
  NOR4_X1   g424(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n601), .A3(new_n602), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n612), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n426), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n276), .A3(new_n436), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n435), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n436), .B1(new_n425), .B2(new_n431), .ZN(new_n621));
  INV_X1    g435(.A(new_n619), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT96), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n392), .A2(new_n570), .A3(new_n598), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT37), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G110), .ZN(G12));
  INV_X1    g442(.A(new_n578), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n574), .A2(new_n188), .A3(new_n575), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n387), .B1(G900), .B2(new_n389), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n507), .A2(new_n521), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n570), .A2(new_n637), .A3(new_n625), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n629), .A2(KEYINPUT97), .A3(new_n630), .A4(new_n633), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XNOR2_X1  g455(.A(new_n631), .B(KEYINPUT98), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT39), .Z(new_n643));
  AND2_X1   g457(.A1(new_n570), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n480), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n492), .B2(new_n516), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n648), .B2(G902), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n507), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n302), .B1(new_n644), .B2(new_n645), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n300), .A2(KEYINPUT38), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n356), .A2(new_n383), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n296), .A2(KEYINPUT38), .A3(new_n299), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n650), .A2(new_n624), .A3(new_n651), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  NOR2_X1   g472(.A1(new_n576), .A2(new_n578), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n589), .B2(new_n631), .ZN(new_n661));
  NOR4_X1   g475(.A1(new_n588), .A2(new_n356), .A3(KEYINPUT99), .A4(new_n632), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(KEYINPUT100), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n629), .A2(new_n630), .A3(new_n663), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n667), .A3(new_n638), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n592), .B2(new_n525), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n276), .B1(new_n552), .B2(new_n555), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(KEYINPUT101), .A3(G469), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n524), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n564), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n671), .A2(new_n673), .B1(new_n558), .B2(new_n563), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n522), .A3(new_n591), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND3_X1  g498(.A1(new_n681), .A2(new_n522), .A3(new_n611), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  INV_X1    g500(.A(new_n676), .ZN(new_n687));
  INV_X1    g501(.A(new_n391), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n624), .B1(new_n507), .B2(new_n521), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n659), .A2(new_n687), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  OAI21_X1  g505(.A(new_n498), .B1(new_n517), .B2(new_n448), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n494), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n597), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n438), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n579), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n576), .A2(new_n578), .A3(new_n654), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n679), .B1(new_n678), .B2(new_n675), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  NOR2_X1   g515(.A1(new_n624), .A2(new_n694), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n659), .A2(new_n687), .A3(new_n663), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  AND3_X1   g518(.A1(new_n296), .A2(new_n301), .A3(new_n299), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n570), .A2(new_n522), .A3(new_n663), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n504), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n438), .B1(new_n709), .B2(new_n521), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n570), .A3(new_n663), .A4(new_n705), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  AND2_X1   g528(.A1(new_n570), .A2(new_n705), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n522), .A3(new_n633), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  XOR2_X1   g531(.A(new_n705), .B(KEYINPUT104), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n585), .A2(new_n587), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n356), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT43), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n624), .A3(new_n598), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n718), .B1(KEYINPUT44), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n567), .B(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(G469), .A2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(G469), .C1(new_n729), .C2(G902), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n564), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(new_n675), .A3(new_n643), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n728), .B(new_n736), .C1(KEYINPUT44), .C2(new_n727), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n675), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n438), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n637), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n663), .A3(new_n705), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  NAND2_X1  g563(.A1(new_n687), .A2(new_n705), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT114), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n507), .A2(new_n649), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n387), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n746), .A3(new_n589), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n384), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT110), .B1(new_n726), .B2(new_n387), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  INV_X1    g571(.A(new_n387), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n724), .A2(new_n757), .A3(new_n758), .A4(new_n725), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n695), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n659), .A3(new_n687), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT118), .Z(new_n762));
  AND3_X1   g576(.A1(new_n755), .A2(KEYINPUT119), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT119), .B1(new_n755), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n759), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n751), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n710), .ZN(new_n767));
  OAI22_X1  g581(.A1(new_n763), .A2(new_n764), .B1(KEYINPUT48), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n687), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n302), .B1(new_n652), .B2(new_n655), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n687), .A4(new_n760), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT113), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n687), .A4(new_n760), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n775), .A3(new_n779), .A4(new_n773), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n766), .A2(new_n702), .ZN(new_n782));
  INV_X1    g596(.A(new_n356), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n719), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n751), .A2(new_n746), .A3(new_n753), .A4(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n781), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  INV_X1    g601(.A(new_n678), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n675), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n745), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n695), .B(new_n718), .C1(new_n759), .C2(new_n756), .ZN(new_n791));
  INV_X1    g605(.A(new_n789), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT116), .B(new_n792), .C1(new_n742), .C2(new_n744), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n786), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n782), .A4(new_n785), .ZN(new_n797));
  INV_X1    g611(.A(new_n794), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n768), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n682), .A2(new_n685), .A3(new_n690), .A4(new_n700), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n570), .A2(new_n663), .A3(new_n705), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n802), .A2(new_n711), .B1(new_n706), .B2(new_n707), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n715), .A2(new_n522), .A3(new_n633), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n702), .A2(new_n570), .A3(new_n663), .A4(new_n705), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n705), .A2(new_n609), .A3(new_n607), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n638), .A2(new_n810), .A3(new_n383), .A4(new_n631), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n801), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n300), .A2(new_n302), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n783), .A2(new_n383), .A3(new_n579), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n601), .A2(new_n814), .A3(new_n602), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n813), .B1(new_n816), .B2(new_n626), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n601), .A2(new_n814), .A3(new_n390), .A4(new_n602), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(new_n590), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n813), .A3(new_n626), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n818), .A2(new_n820), .A3(new_n571), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT109), .B1(new_n812), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n682), .A2(new_n685), .A3(new_n690), .A4(new_n700), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n802), .A2(KEYINPUT108), .A3(new_n702), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n713), .A2(new_n716), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n809), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n816), .A2(new_n813), .A3(new_n626), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n571), .B1(new_n819), .B2(new_n590), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n830), .A3(new_n817), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n831), .A3(new_n832), .A4(new_n811), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n570), .A2(new_n631), .A3(new_n752), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n435), .A3(new_n619), .A4(new_n697), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n668), .A2(new_n640), .A3(new_n835), .A4(new_n703), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n823), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n838), .A2(KEYINPUT53), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n823), .A3(new_n833), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n767), .A2(KEYINPUT48), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n812), .A2(new_n822), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n839), .A2(new_n840), .B1(new_n847), .B2(new_n842), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n800), .A2(new_n845), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n745), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT111), .B1(new_n742), .B2(new_n744), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n792), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n791), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT51), .B1(new_n786), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n851), .A2(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT49), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n596), .B1(new_n678), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n302), .A3(new_n720), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT106), .Z(new_n864));
  NOR2_X1   g678(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n752), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n655), .C2(new_n652), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n210), .A2(G952), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT121), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n842), .A2(new_n847), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n276), .B1(new_n841), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n873), .B2(G210), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n212), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n871), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n841), .A2(new_n872), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(G902), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT120), .B1(new_n848), .B2(new_n276), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n188), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n878), .B1(new_n883), .B2(new_n885), .ZN(G51));
  OR2_X1    g700(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n848), .A2(new_n849), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n841), .A2(new_n849), .A3(new_n872), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n562), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n881), .A2(new_n882), .A3(G469), .A4(new_n729), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n869), .B1(new_n892), .B2(new_n893), .ZN(G54));
  AND2_X1   g708(.A1(KEYINPUT58), .A2(G475), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n881), .A2(new_n882), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n351), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n869), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n881), .A2(new_n882), .A3(new_n351), .A4(new_n895), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G60));
  NAND2_X1  g715(.A1(new_n583), .A2(new_n584), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n380), .A2(new_n276), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n904), .B(new_n905), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n903), .B(new_n907), .C1(new_n889), .C2(new_n890), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n845), .B2(new_n850), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n908), .B(new_n871), .C1(new_n909), .C2(new_n903), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT60), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n879), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n424), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n870), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n841), .B2(new_n872), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n618), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(KEYINPUT124), .A3(new_n618), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n921), .A3(KEYINPUT61), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n871), .B1(new_n918), .B2(new_n424), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT124), .B1(new_n918), .B2(new_n618), .ZN(new_n925));
  INV_X1    g739(.A(new_n618), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n848), .A2(new_n920), .A3(new_n926), .A4(new_n913), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(G66));
  AOI21_X1  g744(.A(new_n210), .B1(new_n388), .B2(G224), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n831), .A2(new_n801), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n875), .B1(G898), .B2(new_n210), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(G69));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n474), .A2(new_n476), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n339), .A2(new_n340), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n668), .A2(new_n640), .A3(new_n703), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n657), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n748), .A2(new_n737), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n590), .B1(new_n383), .B2(new_n783), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n644), .B1(KEYINPUT125), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n946), .A2(new_n522), .A3(new_n705), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n942), .A2(new_n943), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n939), .B1(new_n950), .B2(G953), .ZN(new_n951));
  INV_X1    g765(.A(new_n939), .ZN(new_n952));
  NAND2_X1  g766(.A1(G900), .A2(G953), .ZN(new_n953));
  INV_X1    g767(.A(new_n943), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n803), .A2(new_n804), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n736), .A2(new_n697), .A3(new_n710), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n954), .A2(new_n940), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n952), .B(new_n953), .C1(new_n957), .C2(G953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n936), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n548), .B1(new_n939), .B2(KEYINPUT126), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n210), .B1(new_n960), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  XOR2_X1   g778(.A(new_n941), .B(KEYINPUT62), .Z(new_n965));
  INV_X1    g779(.A(new_n949), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n954), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n967), .B2(new_n932), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n448), .A3(new_n510), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n957), .B2(new_n932), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n492), .A3(new_n509), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n899), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n511), .B(KEYINPUT127), .Z(new_n973));
  AOI22_X1  g787(.A1(new_n841), .A2(new_n843), .B1(new_n480), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n964), .B2(new_n974), .ZN(G57));
endmodule


