

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  AND2_X1 U560 ( .A1(n790), .A2(n1024), .ZN(n526) );
  XOR2_X1 U561 ( .A(n747), .B(KEYINPUT28), .Z(n527) );
  OR2_X1 U562 ( .A1(n794), .A2(n798), .ZN(n528) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n729) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n749) );
  INV_X1 U565 ( .A(KEYINPUT93), .ZN(n765) );
  BUF_X1 U566 ( .A(n755), .Z(n767) );
  INV_X1 U567 ( .A(n798), .ZN(n790) );
  INV_X1 U568 ( .A(KEYINPUT94), .ZN(n784) );
  AND2_X1 U569 ( .A1(n1007), .A2(n528), .ZN(n795) );
  XNOR2_X1 U570 ( .A(n598), .B(KEYINPUT73), .ZN(n736) );
  INV_X1 U571 ( .A(n736), .ZN(n599) );
  NOR2_X2 U572 ( .A1(G651), .A2(n650), .ZN(n658) );
  NOR2_X1 U573 ( .A1(n587), .A2(n586), .ZN(n588) );
  AND2_X1 U574 ( .A1(n545), .A2(n544), .ZN(n690) );
  INV_X1 U575 ( .A(KEYINPUT17), .ZN(n529) );
  XNOR2_X2 U576 ( .A(n530), .B(n529), .ZN(n881) );
  NAND2_X1 U577 ( .A1(G138), .A2(n881), .ZN(n533) );
  INV_X1 U578 ( .A(G2104), .ZN(n531) );
  NOR2_X4 U579 ( .A1(G2105), .A2(n531), .ZN(n882) );
  NAND2_X1 U580 ( .A1(G102), .A2(n882), .ZN(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n538) );
  INV_X1 U582 ( .A(G2105), .ZN(n534) );
  NOR2_X2 U583 ( .A1(n531), .A2(n534), .ZN(n886) );
  NAND2_X1 U584 ( .A1(G114), .A2(n886), .ZN(n536) );
  NOR2_X2 U585 ( .A1(G2104), .A2(n534), .ZN(n887) );
  NAND2_X1 U586 ( .A1(G126), .A2(n887), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U588 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U589 ( .A1(G113), .A2(n886), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G125), .A2(n887), .ZN(n539) );
  AND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n688) );
  NAND2_X1 U592 ( .A1(n881), .A2(G137), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT66), .ZN(n545) );
  NAND2_X1 U594 ( .A1(G101), .A2(n882), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n542), .B(KEYINPUT23), .ZN(n543) );
  XNOR2_X1 U596 ( .A(KEYINPUT65), .B(n543), .ZN(n544) );
  AND2_X1 U597 ( .A1(n688), .A2(n690), .ZN(G160) );
  INV_X1 U598 ( .A(G651), .ZN(n550) );
  NOR2_X1 U599 ( .A1(G543), .A2(n550), .ZN(n547) );
  XNOR2_X1 U600 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n546) );
  XNOR2_X2 U601 ( .A(n547), .B(n546), .ZN(n654) );
  NAND2_X1 U602 ( .A1(G64), .A2(n654), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  NAND2_X1 U604 ( .A1(G52), .A2(n658), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n555) );
  NOR2_X2 U606 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U607 ( .A1(G90), .A2(n653), .ZN(n552) );
  NOR2_X2 U608 ( .A1(n650), .A2(n550), .ZN(n657) );
  NAND2_X1 U609 ( .A1(G77), .A2(n657), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(G62), .A2(n654), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G50), .A2(n658), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT84), .B(n558), .Z(n562) );
  NAND2_X1 U621 ( .A1(G88), .A2(n653), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G75), .A2(n657), .ZN(n559) );
  AND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(G303) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n575) );
  NAND2_X1 U626 ( .A1(n653), .A2(G89), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U628 ( .A1(G76), .A2(n657), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT5), .ZN(n573) );
  XNOR2_X1 U631 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n654), .A2(G63), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT74), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G51), .A2(n658), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n575), .B(n574), .ZN(G168) );
  XOR2_X1 U639 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n577) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G223) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n579) );
  INV_X1 U643 ( .A(G223), .ZN(n831) );
  NAND2_X1 U644 ( .A1(G567), .A2(n831), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G234) );
  NAND2_X1 U646 ( .A1(G68), .A2(n657), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n653), .A2(G81), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G56), .A2(n654), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT14), .B(n584), .Z(n587) );
  NAND2_X1 U653 ( .A1(G43), .A2(n658), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT71), .B(n585), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n1011) );
  INV_X1 U656 ( .A(G860), .ZN(n611) );
  OR2_X1 U657 ( .A1(n1011), .A2(n611), .ZN(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G66), .A2(n654), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G92), .A2(n653), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G79), .A2(n657), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n658), .A2(G54), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT15), .ZN(n598) );
  OR2_X1 U669 ( .A1(n599), .A2(G868), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G284) );
  XOR2_X1 U671 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U672 ( .A1(G65), .A2(n654), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G53), .A2(n658), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G91), .A2(n653), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G78), .A2(n657), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n1015) );
  INV_X1 U679 ( .A(n1015), .ZN(G299) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(G868), .ZN(n608) );
  NOR2_X1 U681 ( .A1(G286), .A2(n608), .ZN(n610) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n612), .A2(n599), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n1011), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G868), .A2(n599), .ZN(n614) );
  NOR2_X1 U689 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U690 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G135), .A2(n881), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G111), .A2(n886), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n887), .A2(G123), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT18), .B(n619), .Z(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n882), .A2(G99), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n976) );
  XOR2_X1 U699 ( .A(G2096), .B(KEYINPUT78), .Z(n624) );
  XNOR2_X1 U700 ( .A(n976), .B(n624), .ZN(n626) );
  INV_X1 U701 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U703 ( .A1(G559), .A2(n599), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(n1011), .ZN(n670) );
  XOR2_X1 U705 ( .A(n670), .B(KEYINPUT79), .Z(n628) );
  NOR2_X1 U706 ( .A1(G860), .A2(n628), .ZN(n629) );
  XOR2_X1 U707 ( .A(KEYINPUT80), .B(n629), .Z(n630) );
  XNOR2_X1 U708 ( .A(KEYINPUT82), .B(n630), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G93), .A2(n653), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G80), .A2(n657), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G67), .A2(n654), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G55), .A2(n658), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U715 ( .A(KEYINPUT81), .B(n635), .Z(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n673) );
  XOR2_X1 U717 ( .A(n638), .B(n673), .Z(G145) );
  NAND2_X1 U718 ( .A1(G86), .A2(n653), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G61), .A2(n654), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n657), .A2(G73), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U724 ( .A(KEYINPUT83), .B(n644), .Z(n646) );
  NAND2_X1 U725 ( .A1(n658), .A2(G48), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n658), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U730 ( .A1(n654), .A2(n649), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(G288) );
  INV_X1 U733 ( .A(G303), .ZN(G166) );
  NAND2_X1 U734 ( .A1(G85), .A2(n653), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G60), .A2(n654), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n662) );
  NAND2_X1 U737 ( .A1(G72), .A2(n657), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G47), .A2(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT68), .B(n663), .Z(G290) );
  XOR2_X1 U742 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n664) );
  XNOR2_X1 U743 ( .A(G288), .B(n664), .ZN(n665) );
  XOR2_X1 U744 ( .A(n665), .B(G166), .Z(n667) );
  XNOR2_X1 U745 ( .A(G290), .B(n1015), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U747 ( .A(n673), .B(n668), .Z(n669) );
  XNOR2_X1 U748 ( .A(G305), .B(n669), .ZN(n902) );
  XNOR2_X1 U749 ( .A(n902), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G868), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(KEYINPUT86), .ZN(n675) );
  OR2_X1 U752 ( .A1(G868), .A2(n673), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2084), .A2(G2078), .ZN(n676) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U762 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G96), .A2(n682), .ZN(n835) );
  NAND2_X1 U764 ( .A1(n835), .A2(G2106), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U766 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G108), .A2(n684), .ZN(n836) );
  NAND2_X1 U768 ( .A1(n836), .A2(G567), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n837) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n837), .A2(n687), .ZN(n834) );
  NAND2_X1 U772 ( .A1(n834), .A2(G36), .ZN(G176) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n722) );
  AND2_X1 U774 ( .A1(n688), .A2(G40), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n722), .A2(n720), .ZN(n826) );
  XNOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  XNOR2_X1 U778 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n886), .A2(G116), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n691), .B(KEYINPUT88), .ZN(n693) );
  NAND2_X1 U781 ( .A1(G128), .A2(n887), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U783 ( .A(n695), .B(n694), .ZN(n701) );
  NAND2_X1 U784 ( .A1(G140), .A2(n881), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G104), .A2(n882), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U787 ( .A(KEYINPUT87), .B(n698), .Z(n699) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n699), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U790 ( .A(KEYINPUT36), .B(n702), .ZN(n898) );
  NOR2_X1 U791 ( .A1(n824), .A2(n898), .ZN(n984) );
  NAND2_X1 U792 ( .A1(n826), .A2(n984), .ZN(n822) );
  NAND2_X1 U793 ( .A1(G131), .A2(n881), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G107), .A2(n886), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U796 ( .A1(G95), .A2(n882), .ZN(n706) );
  NAND2_X1 U797 ( .A1(G119), .A2(n887), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n897) );
  INV_X1 U800 ( .A(G1991), .ZN(n956) );
  NOR2_X1 U801 ( .A1(n897), .A2(n956), .ZN(n717) );
  NAND2_X1 U802 ( .A1(G141), .A2(n881), .ZN(n710) );
  NAND2_X1 U803 ( .A1(G117), .A2(n886), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n882), .A2(G105), .ZN(n711) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n711), .Z(n712) );
  NOR2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n887), .A2(G129), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n878) );
  AND2_X1 U810 ( .A1(G1996), .A2(n878), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n981) );
  INV_X1 U812 ( .A(n826), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n981), .A2(n718), .ZN(n819) );
  INV_X1 U814 ( .A(n819), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n822), .A2(n719), .ZN(n814) );
  INV_X1 U816 ( .A(n720), .ZN(n721) );
  NAND2_X2 U817 ( .A1(n722), .A2(n721), .ZN(n755) );
  AND2_X1 U818 ( .A1(n755), .A2(G1341), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n723), .A2(n1011), .ZN(n728) );
  INV_X1 U820 ( .A(G1996), .ZN(n724) );
  NOR2_X2 U821 ( .A1(n755), .A2(n724), .ZN(n726) );
  XOR2_X1 U822 ( .A(KEYINPUT26), .B(KEYINPUT90), .Z(n725) );
  XNOR2_X1 U823 ( .A(n726), .B(n725), .ZN(n727) );
  AND2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U825 ( .A(n730), .B(n729), .ZN(n737) );
  OR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n735) );
  INV_X1 U827 ( .A(n755), .ZN(n740) );
  INV_X1 U828 ( .A(G1348), .ZN(n1012) );
  NOR2_X1 U829 ( .A1(n740), .A2(n1012), .ZN(n731) );
  XNOR2_X1 U830 ( .A(n731), .B(KEYINPUT91), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n740), .A2(G2067), .ZN(n732) );
  NAND2_X1 U832 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n740), .A2(G2072), .ZN(n741) );
  XNOR2_X1 U837 ( .A(n741), .B(KEYINPUT27), .ZN(n743) );
  AND2_X1 U838 ( .A1(G1956), .A2(n767), .ZN(n742) );
  NOR2_X1 U839 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n1015), .A2(n746), .ZN(n744) );
  NAND2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n1015), .A2(n746), .ZN(n747) );
  NAND2_X1 U843 ( .A1(n748), .A2(n527), .ZN(n750) );
  XNOR2_X1 U844 ( .A(n750), .B(n749), .ZN(n754) );
  INV_X1 U845 ( .A(G1961), .ZN(n925) );
  NAND2_X1 U846 ( .A1(n767), .A2(n925), .ZN(n752) );
  XNOR2_X1 U847 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U848 ( .A1(n740), .A2(n955), .ZN(n751) );
  NAND2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n759), .A2(G171), .ZN(n753) );
  NAND2_X1 U851 ( .A1(n754), .A2(n753), .ZN(n764) );
  NOR2_X1 U852 ( .A1(G2084), .A2(n767), .ZN(n779) );
  NAND2_X1 U853 ( .A1(G8), .A2(n755), .ZN(n798) );
  NOR2_X1 U854 ( .A1(G1966), .A2(n798), .ZN(n777) );
  NOR2_X1 U855 ( .A1(n779), .A2(n777), .ZN(n756) );
  NAND2_X1 U856 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U857 ( .A(KEYINPUT30), .B(n757), .ZN(n758) );
  NOR2_X1 U858 ( .A1(G168), .A2(n758), .ZN(n761) );
  NOR2_X1 U859 ( .A1(G171), .A2(n759), .ZN(n760) );
  NOR2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U861 ( .A(KEYINPUT31), .B(n762), .Z(n763) );
  NAND2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n775), .A2(G286), .ZN(n766) );
  XNOR2_X1 U864 ( .A(n766), .B(n765), .ZN(n772) );
  NOR2_X1 U865 ( .A1(G1971), .A2(n798), .ZN(n769) );
  NOR2_X1 U866 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U867 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U868 ( .A1(G303), .A2(n770), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n773), .A2(G8), .ZN(n774) );
  XNOR2_X1 U871 ( .A(n774), .B(KEYINPUT32), .ZN(n783) );
  INV_X1 U872 ( .A(n775), .ZN(n776) );
  NOR2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U874 ( .A(n778), .B(KEYINPUT92), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n779), .A2(G8), .ZN(n780) );
  NAND2_X1 U876 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n785) );
  XNOR2_X2 U878 ( .A(n785), .B(n784), .ZN(n802) );
  NOR2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n1022) );
  NOR2_X2 U880 ( .A1(n802), .A2(n1022), .ZN(n788) );
  NOR2_X1 U881 ( .A1(G1971), .A2(G303), .ZN(n786) );
  XNOR2_X1 U882 ( .A(n786), .B(KEYINPUT95), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G288), .A2(G1976), .ZN(n789) );
  XNOR2_X1 U885 ( .A(n789), .B(KEYINPUT96), .ZN(n1024) );
  NAND2_X1 U886 ( .A1(n791), .A2(n526), .ZN(n793) );
  INV_X1 U887 ( .A(KEYINPUT33), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n796) );
  XOR2_X1 U889 ( .A(G1981), .B(G305), .Z(n1007) );
  NAND2_X1 U890 ( .A1(n1022), .A2(KEYINPUT33), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U892 ( .A(n797), .B(KEYINPUT97), .ZN(n811) );
  INV_X1 U893 ( .A(G8), .ZN(n801) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n799) );
  XOR2_X1 U895 ( .A(KEYINPUT98), .B(n799), .Z(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n790), .A2(n804), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(KEYINPUT99), .ZN(n809) );
  NOR2_X1 U900 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT24), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n790), .A2(n807), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT100), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U907 ( .A(G290), .B(G1986), .ZN(n1014) );
  NAND2_X1 U908 ( .A1(n1014), .A2(n826), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n829) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n878), .ZN(n987) );
  NOR2_X1 U911 ( .A1(G290), .A2(G1986), .ZN(n817) );
  AND2_X1 U912 ( .A1(n956), .A2(n897), .ZN(n979) );
  NOR2_X1 U913 ( .A1(n817), .A2(n979), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n987), .A2(n820), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n824), .A2(n898), .ZN(n992) );
  NAND2_X1 U919 ( .A1(n825), .A2(n992), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n837), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT41), .B(G1966), .Z(n839) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n840), .B(KEYINPUT106), .Z(n842) );
  XNOR2_X1 U939 ( .A(G1956), .B(G1976), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(G1971), .B(G1961), .Z(n844) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1981), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(G2474), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2100), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(KEYINPUT103), .B(G2090), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT104), .B(G2096), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U956 ( .A(G2084), .B(G2078), .Z(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G100), .A2(n882), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G112), .A2(n886), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n887), .A2(G124), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G136), .A2(n881), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(KEYINPUT107), .B(n864), .Z(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n877) );
  NAND2_X1 U968 ( .A1(G118), .A2(n886), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G130), .A2(n887), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G142), .A2(n881), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G106), .A2(n882), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(KEYINPUT108), .B(n871), .Z(n872) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n872), .ZN(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n896) );
  XOR2_X1 U979 ( .A(G160), .B(n878), .Z(n879) );
  XNOR2_X1 U980 ( .A(n879), .B(G162), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n976), .B(n880), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G139), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT109), .B(n885), .Z(n892) );
  NAND2_X1 U986 ( .A1(G115), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G127), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n994) );
  XNOR2_X1 U991 ( .A(G164), .B(n994), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U997 ( .A(n1011), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(G171), .B(n599), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(G286), .Z(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U1002 ( .A(G2451), .B(G2446), .ZN(n916) );
  XOR2_X1 U1003 ( .A(G2430), .B(G2443), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2435), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1006 ( .A(G2438), .B(KEYINPUT101), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT102), .B(G2427), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n917), .A2(G14), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT111), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n924), .ZN(G401) );
  XNOR2_X1 U1024 ( .A(G5), .B(n925), .ZN(n946) );
  XNOR2_X1 U1025 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n936) );
  XNOR2_X1 U1026 ( .A(KEYINPUT59), .B(G1348), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n926), .B(G4), .ZN(n934) );
  XOR2_X1 U1028 ( .A(G1341), .B(G19), .Z(n929) );
  XOR2_X1 U1029 ( .A(G20), .B(KEYINPUT124), .Z(n927) );
  XNOR2_X1 U1030 ( .A(G1956), .B(n927), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1032 ( .A(KEYINPUT125), .B(G1981), .Z(n930) );
  XNOR2_X1 U1033 ( .A(G6), .B(n930), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G1986), .B(G24), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G22), .B(G1971), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G1976), .B(KEYINPUT127), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(n939), .B(G23), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(n942), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G21), .B(G1966), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1048 ( .A(KEYINPUT61), .B(n949), .Z(n950) );
  NOR2_X1 U1049 ( .A1(G16), .A2(n950), .ZN(n975) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1002) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n951), .ZN(n968) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n966) );
  XOR2_X1 U1054 ( .A(G2067), .B(G26), .Z(n952) );
  NAND2_X1 U1055 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1057 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1058 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1059 ( .A(n955), .B(G27), .Z(n958) );
  XOR2_X1 U1060 ( .A(n956), .B(G25), .Z(n957) );
  NOR2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1062 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1064 ( .A(KEYINPUT53), .B(n963), .Z(n964) );
  XNOR2_X1 U1065 ( .A(n964), .B(KEYINPUT117), .ZN(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(n1002), .B(n969), .ZN(n970) );
  XNOR2_X1 U1069 ( .A(KEYINPUT118), .B(n970), .ZN(n972) );
  INV_X1 U1070 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1072 ( .A1(n973), .A2(G11), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n1006) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n977) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT112), .B(n980), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT113), .B(n985), .ZN(n990) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(KEYINPUT51), .B(n988), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n991), .B(KEYINPUT114), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G2072), .B(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G164), .B(G2078), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT115), .B(n997), .Z(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT50), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(G29), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1038) );
  XOR2_X1 U1097 ( .A(KEYINPUT56), .B(G16), .Z(n1036) );
  XNOR2_X1 U1098 ( .A(KEYINPUT57), .B(KEYINPUT119), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1010), .B(n1009), .ZN(n1033) );
  XNOR2_X1 U1102 ( .A(n1011), .B(G1341), .ZN(n1030) );
  XNOR2_X1 U1103 ( .A(n599), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1015), .B(G1956), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G171), .B(G1961), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(G1971), .B(G303), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1027) );
  INV_X1 U1111 ( .A(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT120), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT121), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT122), .B(n1031), .Z(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT123), .B(n1034), .Z(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1122 ( .A(n1039), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

