//key=1010101010101010101010101010101010101010101010101010101010101010


module locked_locked_c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, 
        G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, 
        G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, 
        G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, 
        G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, 
        G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, 
        G409, G405, G402, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, 
        KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, 
        KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, 
        KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, 
        KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, 
        KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, 
        KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, 
        KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, 
        KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, 
        KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, 
        KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, 
        KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, 
        KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, 
        KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, 
        KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, 
        KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, 
        KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, 
        KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, 
        KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, 
        KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, 
        KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, 
        KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, 
        KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60,
         KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55,
         KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50,
         KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45,
         KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40,
         KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35,
         KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30,
         KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25,
         KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20,
         KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15,
         KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9,
         KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3,
         KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126,
         KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121,
         KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116,
         KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111,
         KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106,
         KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101,
         KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96,
         KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91,
         KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86,
         KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81,
         KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76,
         KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71,
         KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66,
         KEYINPUT65, KEYINPUT64;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
         G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071;

  NOR2_X1 U1034 ( .A1(n1133), .A2(n1132), .ZN(n1136) );
  NAND2_X1 U1035 ( .A1(n1525), .A2(n1524), .ZN(n1674) );
  NAND2_X1 U1036 ( .A1(n1078), .A2(n1033), .ZN(G378) );
  INV_X1 U1037 ( .A(n2071), .ZN(n1063) );
  NOR2_X2 U1038 ( .A1(n1484), .A2(n1542), .ZN(n1522) );
  NAND2_X2 U1039 ( .A1(G13), .A2(G1), .ZN(n1103) );
  NAND2_X1 U1040 ( .A1(n1079), .A2(n1605), .ZN(G375) );
  AND2_X2 U1041 ( .A1(n1521), .A2(n1416), .ZN(n1542) );
  NOR2_X2 U1042 ( .A1(n1123), .A2(n1122), .ZN(n1239) );
  XNOR2_X2 U1043 ( .A(n1232), .B(KEYINPUT77), .ZN(n1259) );
  OR2_X1 U1044 ( .A1(n1355), .A2(n1354), .ZN(G390) );
  XNOR2_X1 U1045 ( .A(n1857), .B(KEYINPUT55), .ZN(G387) );
  XNOR2_X1 U1046 ( .A(n1072), .B(n1527), .ZN(n1715) );
  AND2_X1 U1047 ( .A1(n1492), .A2(n1491), .ZN(n2018) );
  OR2_X2 U1048 ( .A1(n1209), .A2(n1246), .ZN(n1293) );
  NOR2_X1 U1049 ( .A1(n1140), .A2(n1137), .ZN(n1040) );
  OR2_X1 U1050 ( .A1(n1259), .A2(n1084), .ZN(n1234) );
  XNOR2_X1 U1051 ( .A(n1088), .B(KEYINPUT69), .ZN(n1372) );
  AND2_X1 U1052 ( .A1(n1991), .A2(n1044), .ZN(n1023) );
  INV_X1 U1053 ( .A(n1119), .ZN(n1991) );
  NAND2_X1 U1054 ( .A1(n1163), .A2(n1162), .ZN(n1180) );
  NAND2_X1 U1055 ( .A1(n1164), .A2(n1180), .ZN(n1211) );
  XNOR2_X1 U1056 ( .A(n1261), .B(n1038), .ZN(n1262) );
  INV_X1 U1057 ( .A(KEYINPUT18), .ZN(n1038) );
  NOR2_X1 U1058 ( .A1(n1260), .A2(n1259), .ZN(n1261) );
  NAND2_X1 U1059 ( .A1(n1068), .A2(n1031), .ZN(n1503) );
  INV_X1 U1060 ( .A(n1500), .ZN(n1068) );
  NAND2_X1 U1061 ( .A1(n1024), .A2(n1015), .ZN(n1494) );
  AND2_X1 U1062 ( .A1(n1283), .A2(n1669), .ZN(n1218) );
  AND2_X1 U1063 ( .A1(n1090), .A2(n1018), .ZN(n1216) );
  NAND2_X1 U1064 ( .A1(n1266), .A2(n1021), .ZN(n1090) );
  NAND2_X1 U1065 ( .A1(n1021), .A2(n1184), .ZN(n1089) );
  OR2_X1 U1066 ( .A1(n1253), .A2(n1784), .ZN(n1495) );
  AND2_X1 U1067 ( .A1(n1388), .A2(n1387), .ZN(n1556) );
  NAND2_X1 U1068 ( .A1(n1991), .A2(n1110), .ZN(n1088) );
  NAND2_X1 U1069 ( .A1(n1037), .A2(n2043), .ZN(n1534) );
  NAND2_X1 U1070 ( .A1(n1016), .A2(n1025), .ZN(n1037) );
  NAND2_X1 U1071 ( .A1(n2016), .A2(n1796), .ZN(n1533) );
  NOR2_X1 U1072 ( .A1(n1047), .A2(n1046), .ZN(n1049) );
  OR2_X1 U1073 ( .A1(n1019), .A2(G179), .ZN(n1046) );
  NAND2_X1 U1074 ( .A1(n1045), .A2(n1020), .ZN(n1264) );
  NOR2_X1 U1075 ( .A1(n1109), .A2(n1019), .ZN(n1045) );
  NOR2_X1 U1076 ( .A1(n1152), .A2(n1151), .ZN(n1154) );
  NOR2_X1 U1077 ( .A1(n1507), .A2(n1506), .ZN(n1540) );
  INV_X1 U1078 ( .A(n1494), .ZN(n1501) );
  XNOR2_X1 U1079 ( .A(n1144), .B(n1143), .ZN(n1214) );
  XNOR2_X1 U1080 ( .A(n1142), .B(KEYINPUT66), .ZN(n1143) );
  OR2_X1 U1081 ( .A1(n1512), .A2(n1508), .ZN(n1498) );
  XNOR2_X1 U1082 ( .A(n1041), .B(G396), .ZN(n1054) );
  XNOR2_X1 U1083 ( .A(n1210), .B(n1293), .ZN(n1283) );
  OR2_X1 U1084 ( .A1(n1219), .A2(n1293), .ZN(n1786) );
  XNOR2_X1 U1085 ( .A(n1252), .B(KEYINPUT67), .ZN(n1784) );
  XNOR2_X1 U1086 ( .A(n1183), .B(KEYINPUT11), .ZN(n1266) );
  NOR2_X1 U1087 ( .A1(n1182), .A2(n1181), .ZN(n1183) );
  NAND2_X1 U1088 ( .A1(n1498), .A2(n1496), .ZN(n1510) );
  NAND2_X1 U1089 ( .A1(n1477), .A2(n1494), .ZN(n1500) );
  NOR2_X1 U1090 ( .A1(n1389), .A2(n1556), .ZN(n1390) );
  NAND2_X1 U1091 ( .A1(n1063), .A2(n1036), .ZN(n1060) );
  NAND2_X1 U1092 ( .A1(n1059), .A2(n1057), .ZN(n1056) );
  NAND2_X1 U1093 ( .A1(n1916), .A2(KEYINPUT125), .ZN(n1059) );
  NAND2_X1 U1094 ( .A1(n1066), .A2(n1058), .ZN(n1057) );
  NAND2_X1 U1095 ( .A1(n1914), .A2(KEYINPUT125), .ZN(n1058) );
  XNOR2_X1 U1096 ( .A(n1061), .B(n1064), .ZN(n2070) );
  XNOR2_X1 U1097 ( .A(G381), .B(G393), .ZN(n1064) );
  XNOR2_X1 U1098 ( .A(G387), .B(n1053), .ZN(n1061) );
  XNOR2_X1 U1099 ( .A(G390), .B(n1054), .ZN(n1053) );
  AND2_X1 U1100 ( .A1(n1560), .A2(n1940), .ZN(n1080) );
  NOR2_X1 U1101 ( .A1(n1096), .A2(n2023), .ZN(n1093) );
  INV_X1 U1102 ( .A(G270), .ZN(n1087) );
  AND2_X1 U1103 ( .A1(n1991), .A2(n1042), .ZN(n1145) );
  AND2_X1 U1104 ( .A1(n1043), .A2(G33), .ZN(n1042) );
  INV_X1 U1105 ( .A(G41), .ZN(n1043) );
  AND2_X1 U1106 ( .A1(n1120), .A2(n1289), .ZN(n1129) );
  XNOR2_X1 U1107 ( .A(n1118), .B(n1117), .ZN(n1120) );
  BUF_X2 U1108 ( .A(n1445), .Z(n1434) );
  INV_X1 U1109 ( .A(KEYINPUT65), .ZN(n1052) );
  NAND2_X1 U1110 ( .A1(n1495), .A2(n1077), .ZN(n1074) );
  AND2_X1 U1111 ( .A1(n1496), .A2(n1796), .ZN(n1077) );
  AND2_X1 U1112 ( .A1(n1121), .A2(G33), .ZN(n1044) );
  INV_X1 U1113 ( .A(KEYINPUT36), .ZN(n1377) );
  NOR2_X1 U1114 ( .A1(n1375), .A2(n1374), .ZN(n1376) );
  NOR2_X1 U1115 ( .A1(n1231), .A2(n1230), .ZN(n1232) );
  OR2_X1 U1116 ( .A1(n1393), .A2(n1239), .ZN(n1156) );
  NAND2_X1 U1117 ( .A1(n1075), .A2(n1073), .ZN(n1529) );
  NAND2_X1 U1118 ( .A1(n1786), .A2(n1076), .ZN(n1075) );
  NAND2_X1 U1119 ( .A1(n1074), .A2(n1499), .ZN(n1073) );
  AND2_X1 U1120 ( .A1(n1499), .A2(n1247), .ZN(n1076) );
  AND2_X1 U1121 ( .A1(n1503), .A2(n1502), .ZN(n1505) );
  AND2_X1 U1122 ( .A1(n1153), .A2(G179), .ZN(n1082) );
  NAND2_X1 U1123 ( .A1(n1269), .A2(n1533), .ZN(n1528) );
  XNOR2_X1 U1124 ( .A(n1049), .B(KEYINPUT15), .ZN(n1139) );
  XNOR2_X1 U1125 ( .A(n1382), .B(n1381), .ZN(n1386) );
  INV_X1 U1126 ( .A(KEYINPUT99), .ZN(n1381) );
  NOR2_X1 U1127 ( .A1(n1380), .A2(n1379), .ZN(n1382) );
  XNOR2_X1 U1128 ( .A(n1378), .B(n1377), .ZN(n1379) );
  NAND2_X1 U1129 ( .A1(n1202), .A2(n1201), .ZN(n1260) );
  XNOR2_X1 U1130 ( .A(KEYINPUT12), .B(KEYINPUT74), .ZN(n1198) );
  XNOR2_X1 U1131 ( .A(n1674), .B(n1526), .ZN(n1527) );
  INV_X1 U1132 ( .A(n2026), .ZN(n1096) );
  OR2_X1 U1133 ( .A1(n1912), .A2(n1911), .ZN(n1041) );
  OR2_X1 U1134 ( .A1(n1266), .A2(n1184), .ZN(n1091) );
  AND2_X1 U1135 ( .A1(n1497), .A2(n1495), .ZN(n1050) );
  NOR2_X1 U1136 ( .A1(n1482), .A2(n1556), .ZN(n2042) );
  INV_X1 U1137 ( .A(n1214), .ZN(n1268) );
  INV_X1 U1138 ( .A(n1510), .ZN(n1490) );
  AND2_X1 U1139 ( .A1(G1), .A2(G20), .ZN(n1101) );
  NAND2_X1 U1140 ( .A1(n2071), .A2(n1035), .ZN(n1055) );
  NAND2_X1 U1141 ( .A1(n1081), .A2(n1080), .ZN(n1079) );
  AND2_X1 U1142 ( .A1(n1278), .A2(n1097), .ZN(n1355) );
  NOR2_X1 U1143 ( .A1(n1667), .A2(n1666), .ZN(n1668) );
  NOR2_X1 U1144 ( .A1(n1856), .A2(n1855), .ZN(n1857) );
  AND2_X1 U1145 ( .A1(n1095), .A2(n1028), .ZN(n1856) );
  INV_X1 U1146 ( .A(n1041), .ZN(G384) );
  XNOR2_X1 U1147 ( .A(n1505), .B(n1504), .ZN(n1531) );
  OR2_X1 U1148 ( .A1(n1431), .A2(n1430), .ZN(n1015) );
  OR2_X1 U1149 ( .A1(n1265), .A2(n1264), .ZN(n1016) );
  XNOR2_X1 U1150 ( .A(G375), .B(G378), .ZN(n2071) );
  AND2_X1 U1151 ( .A1(n1439), .A2(n1029), .ZN(n1017) );
  AND2_X1 U1152 ( .A1(n1089), .A2(G330), .ZN(n1018) );
  INV_X1 U1153 ( .A(KEYINPUT125), .ZN(n1065) );
  AND2_X1 U1154 ( .A1(n1448), .A2(G257), .ZN(n1019) );
  AND2_X1 U1155 ( .A1(n1192), .A2(n1112), .ZN(n1020) );
  OR2_X1 U1156 ( .A1(n1211), .A2(n1796), .ZN(n1021) );
  AND2_X1 U1157 ( .A1(n1091), .A2(n1021), .ZN(n1022) );
  AND2_X1 U1158 ( .A1(n1443), .A2(n1442), .ZN(n1024) );
  OR2_X1 U1159 ( .A1(n1258), .A2(n1257), .ZN(n1025) );
  OR2_X1 U1160 ( .A1(n1714), .A2(n1713), .ZN(n1026) );
  AND2_X1 U1161 ( .A1(n1386), .A2(n1084), .ZN(n1027) );
  XNOR2_X1 U1162 ( .A(n1802), .B(n1801), .ZN(n1028) );
  AND2_X1 U1163 ( .A1(n1440), .A2(n1084), .ZN(n1029) );
  OR2_X1 U1164 ( .A1(n1260), .A2(n1083), .ZN(n1030) );
  NAND2_X1 U1165 ( .A1(n1015), .A2(n2043), .ZN(n1031) );
  AND2_X1 U1166 ( .A1(n1153), .A2(G190), .ZN(n1032) );
  AND2_X1 U1167 ( .A1(n1719), .A2(n1026), .ZN(n1033) );
  AND2_X1 U1168 ( .A1(n1060), .A2(n1056), .ZN(n1034) );
  INV_X1 U1169 ( .A(G190), .ZN(n1083) );
  NOR2_X1 U1170 ( .A1(n1992), .A2(G41), .ZN(n2031) );
  INV_X1 U1171 ( .A(n1916), .ZN(n1066) );
  AND2_X1 U1172 ( .A1(n1066), .A2(KEYINPUT125), .ZN(n1035) );
  BUF_X1 U1173 ( .A(G1), .Z(n2022) );
  AND2_X1 U1174 ( .A1(n1067), .A2(n1065), .ZN(n1036) );
  NOR2_X2 U1175 ( .A1(n1084), .A2(n1319), .ZN(n1947) );
  NOR2_X2 U1176 ( .A1(n1084), .A2(n1303), .ZN(n1953) );
  NOR2_X2 U1177 ( .A1(G179), .A2(n1319), .ZN(n1946) );
  NOR2_X2 U1178 ( .A1(n1084), .A2(n1302), .ZN(n1952) );
  NOR2_X2 U1179 ( .A1(n1311), .A2(n1297), .ZN(n1956) );
  NOR2_X2 U1180 ( .A1(G179), .A2(n1303), .ZN(n1943) );
  NAND2_X1 U1181 ( .A1(n1039), .A2(n1517), .ZN(n1530) );
  INV_X1 U1182 ( .A(n1528), .ZN(n1039) );
  NAND2_X1 U1183 ( .A1(G407), .A2(n1990), .ZN(G409) );
  NAND2_X1 U1184 ( .A1(n1985), .A2(n1986), .ZN(G407) );
  NOR2_X1 U1185 ( .A1(n1197), .A2(n1196), .ZN(n1199) );
  NAND2_X1 U1186 ( .A1(n1040), .A2(n2043), .ZN(n1186) );
  NOR2_X1 U1187 ( .A1(n1141), .A2(n1040), .ZN(n1144) );
  NOR2_X1 U1188 ( .A1(n1165), .A2(n1040), .ZN(n1219) );
  NOR2_X1 U1189 ( .A1(G387), .A2(G384), .ZN(n1981) );
  NAND2_X1 U1190 ( .A1(n1048), .A2(n1020), .ZN(n1047) );
  INV_X1 U1191 ( .A(n1109), .ZN(n1048) );
  NAND2_X1 U1192 ( .A1(n1050), .A2(n1796), .ZN(n1270) );
  NAND2_X1 U1193 ( .A1(n2018), .A2(n1050), .ZN(n1493) );
  AND2_X2 U1194 ( .A1(n1051), .A2(n1108), .ZN(n1148) );
  AND2_X2 U1195 ( .A1(n1051), .A2(G1698), .ZN(n1448) );
  AND2_X1 U1196 ( .A1(n1051), .A2(n1121), .ZN(n1466) );
  XNOR2_X2 U1197 ( .A(n1105), .B(n1052), .ZN(n1051) );
  NAND2_X1 U1198 ( .A1(n1034), .A2(n1055), .ZN(n1062) );
  XNOR2_X1 U1199 ( .A(n1062), .B(n2070), .ZN(G405) );
  INV_X1 U1200 ( .A(n1914), .ZN(n1067) );
  NAND2_X1 U1201 ( .A1(n1439), .A2(n1440), .ZN(n1069) );
  NAND2_X1 U1202 ( .A1(n1069), .A2(G200), .ZN(n1473) );
  NOR2_X1 U1203 ( .A1(n1069), .A2(n1083), .ZN(n1472) );
  NAND2_X1 U1204 ( .A1(n1069), .A2(n1441), .ZN(n1442) );
  XNOR2_X1 U1205 ( .A(n1071), .B(n1070), .ZN(n1539) );
  INV_X1 U1206 ( .A(KEYINPUT41), .ZN(n1070) );
  NAND2_X1 U1207 ( .A1(n1715), .A2(n1972), .ZN(n1071) );
  NAND2_X1 U1208 ( .A1(n1520), .A2(n1540), .ZN(n1072) );
  NOR2_X2 U1209 ( .A1(n2019), .A2(n1294), .ZN(n1188) );
  NOR2_X1 U1210 ( .A1(G390), .A2(G381), .ZN(n1982) );
  NOR2_X1 U1211 ( .A1(n1920), .A2(n2023), .ZN(n1921) );
  NAND2_X1 U1212 ( .A1(n1795), .A2(n1798), .ZN(n1251) );
  NAND2_X1 U1213 ( .A1(n1786), .A2(n1247), .ZN(n1497) );
  NOR2_X2 U1214 ( .A1(n1413), .A2(n1084), .ZN(n1412) );
  NAND2_X1 U1215 ( .A1(n1718), .A2(n2031), .ZN(n1078) );
  NAND2_X1 U1216 ( .A1(n1539), .A2(n1538), .ZN(n1081) );
  NAND2_X1 U1217 ( .A1(n1154), .A2(n1153), .ZN(n1176) );
  NAND2_X1 U1218 ( .A1(n1154), .A2(n1032), .ZN(n1177) );
  NAND2_X1 U1219 ( .A1(n1154), .A2(n1082), .ZN(n1263) );
  AND2_X1 U1220 ( .A1(n1176), .A2(n1084), .ZN(n1255) );
  INV_X1 U1221 ( .A(G179), .ZN(n1084) );
  XNOR2_X1 U1222 ( .A(n2070), .B(n1063), .ZN(G402) );
  NAND2_X1 U1223 ( .A1(n1085), .A2(n1086), .ZN(n1147) );
  INV_X1 U1224 ( .A(n1372), .ZN(n1085) );
  NOR2_X1 U1225 ( .A1(n1372), .A2(n1111), .ZN(n1200) );
  NOR2_X1 U1226 ( .A1(n1111), .A2(n1087), .ZN(n1086) );
  NAND2_X1 U1227 ( .A1(n1094), .A2(n1092), .ZN(n1095) );
  NOR2_X1 U1228 ( .A1(n1093), .A2(n1973), .ZN(n1092) );
  NAND2_X1 U1229 ( .A1(n1782), .A2(n2031), .ZN(n1094) );
  NOR2_X1 U1230 ( .A1(n1438), .A2(n1437), .ZN(n1439) );
  AND2_X1 U1231 ( .A1(n1522), .A2(n1490), .ZN(n1491) );
  NAND2_X1 U1232 ( .A1(n1100), .A2(n1268), .ZN(n2016) );
  NOR2_X1 U1233 ( .A1(n1518), .A2(n1528), .ZN(n1519) );
  NAND2_X1 U1234 ( .A1(n1270), .A2(n1528), .ZN(n2026) );
  AND2_X1 U1235 ( .A1(n1277), .A2(n2031), .ZN(n1097) );
  OR2_X1 U1236 ( .A1(n1372), .A2(n1228), .ZN(n1098) );
  INV_X1 U1237 ( .A(n1129), .ZN(n1359) );
  OR2_X1 U1238 ( .A1(G116), .A2(n1462), .ZN(n1099) );
  AND2_X1 U1239 ( .A1(n1267), .A2(n1784), .ZN(n1100) );
  INV_X1 U1240 ( .A(KEYINPUT6), .ZN(n1449) );
  INV_X1 U1241 ( .A(KEYINPUT3), .ZN(n1117) );
  INV_X1 U1242 ( .A(G20), .ZN(n1121) );
  AND2_X1 U1243 ( .A1(n1099), .A2(n1158), .ZN(n1159) );
  BUF_X1 U1244 ( .A(n1119), .Z(n1289) );
  NOR2_X1 U1245 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
  INV_X1 U1246 ( .A(KEYINPUT38), .ZN(n1536) );
  INV_X1 U1247 ( .A(KEYINPUT40), .ZN(n1526) );
  INV_X1 U1248 ( .A(KEYINPUT0), .ZN(n1142) );
  INV_X1 U1249 ( .A(G13), .ZN(n1287) );
  NOR2_X1 U1250 ( .A1(G20), .A2(n1287), .ZN(n1279) );
  NAND2_X1 U1251 ( .A1(n1279), .A2(G213), .ZN(n1102) );
  NOR2_X1 U1252 ( .A1(n2022), .A2(n1102), .ZN(n1555) );
  NAND2_X1 U1253 ( .A1(n1555), .A2(G343), .ZN(n1796) );
  INV_X1 U1254 ( .A(n1796), .ZN(n2043) );
  XNOR2_X2 U1255 ( .A(n1103), .B(KEYINPUT2), .ZN(n1119) );
  NAND2_X1 U1256 ( .A1(n1145), .A2(G294), .ZN(n1104) );
  XNOR2_X1 U1257 ( .A(n1104), .B(KEYINPUT14), .ZN(n1107) );
  NOR2_X2 U1258 ( .A1(n1119), .A2(G33), .ZN(n1105) );
  NAND2_X1 U1259 ( .A1(G250), .A2(n1148), .ZN(n1106) );
  NAND2_X1 U1260 ( .A1(n1107), .A2(n1106), .ZN(n1109) );
  INV_X1 U1261 ( .A(G1698), .ZN(n1108) );
  INV_X1 U1262 ( .A(n2022), .ZN(n2027) );
  NAND2_X1 U1263 ( .A1(G45), .A2(n2027), .ZN(n1227) );
  NOR2_X1 U1264 ( .A1(G41), .A2(n1227), .ZN(n1111) );
  NAND2_X1 U1265 ( .A1(G274), .A2(n1111), .ZN(n1192) );
  NAND2_X1 U1266 ( .A1(G33), .A2(G41), .ZN(n1110) );
  NAND2_X1 U1267 ( .A1(G264), .A2(n1200), .ZN(n1112) );
  NOR2_X1 U1268 ( .A1(n1264), .A2(n1083), .ZN(n1113) );
  XNOR2_X1 U1269 ( .A(n1113), .B(KEYINPUT71), .ZN(n1115) );
  NAND2_X1 U1270 ( .A1(n1264), .A2(G200), .ZN(n1114) );
  NAND2_X1 U1271 ( .A1(n1115), .A2(n1114), .ZN(n1135) );
  NAND2_X1 U1272 ( .A1(G116), .A2(n1023), .ZN(n1116) );
  XNOR2_X1 U1273 ( .A(n1116), .B(KEYINPUT16), .ZN(n1125) );
  NAND2_X1 U1274 ( .A1(n1101), .A2(G33), .ZN(n1118) );
  NOR2_X1 U1275 ( .A1(n2022), .A2(n1121), .ZN(n1360) );
  NAND2_X1 U1276 ( .A1(G13), .A2(n1360), .ZN(n1462) );
  NAND2_X1 U1277 ( .A1(n1129), .A2(n1462), .ZN(n1123) );
  INV_X1 U1278 ( .A(G33), .ZN(n1898) );
  NOR2_X1 U1279 ( .A1(n2022), .A2(n1898), .ZN(n1122) );
  NAND2_X1 U1280 ( .A1(n1239), .A2(G107), .ZN(n1124) );
  NAND2_X1 U1281 ( .A1(n1125), .A2(n1124), .ZN(n1126) );
  XNOR2_X1 U1282 ( .A(n1126), .B(KEYINPUT17), .ZN(n1128) );
  NAND2_X1 U1283 ( .A1(n1466), .A2(G87), .ZN(n1127) );
  NAND2_X1 U1284 ( .A1(n1128), .A2(n1127), .ZN(n1133) );
  INV_X1 U1285 ( .A(n1462), .ZN(n1356) );
  NAND2_X1 U1286 ( .A1(G20), .A2(n1359), .ZN(n1131) );
  INV_X1 U1287 ( .A(KEYINPUT4), .ZN(n1130) );
  XNOR2_X2 U1288 ( .A(n1131), .B(n1130), .ZN(n1393) );
  NOR2_X1 U1289 ( .A1(n1356), .A2(n1393), .ZN(n1429) );
  NOR2_X1 U1290 ( .A1(G107), .A2(n1429), .ZN(n1132) );
  XOR2_X1 U1291 ( .A(n1136), .B(KEYINPUT70), .Z(n1134) );
  NOR2_X1 U1292 ( .A1(n1135), .A2(n1134), .ZN(n1141) );
  BUF_X1 U1293 ( .A(n1136), .Z(n1137) );
  INV_X1 U1294 ( .A(G169), .ZN(n1441) );
  NAND2_X1 U1295 ( .A1(n1264), .A2(n1441), .ZN(n1138) );
  NAND2_X1 U1296 ( .A1(n1139), .A2(n1138), .ZN(n1140) );
  XNOR2_X2 U1297 ( .A(n1145), .B(KEYINPUT68), .ZN(n1444) );
  NAND2_X1 U1298 ( .A1(G303), .A2(n1444), .ZN(n1146) );
  NAND2_X1 U1299 ( .A1(n1192), .A2(n1146), .ZN(n1152) );
  XNOR2_X1 U1300 ( .A(n1147), .B(KEYINPUT10), .ZN(n1150) );
  XNOR2_X2 U1301 ( .A(n1148), .B(KEYINPUT64), .ZN(n1445) );
  NAND2_X1 U1302 ( .A1(G257), .A2(n1445), .ZN(n1149) );
  NAND2_X1 U1303 ( .A1(n1150), .A2(n1149), .ZN(n1151) );
  NAND2_X1 U1304 ( .A1(n1448), .A2(G264), .ZN(n1153) );
  NAND2_X1 U1305 ( .A1(n1176), .A2(G169), .ZN(n1155) );
  NAND2_X1 U1306 ( .A1(n1155), .A2(n1263), .ZN(n1164) );
  NAND2_X1 U1307 ( .A1(n1156), .A2(G116), .ZN(n1157) );
  XNOR2_X1 U1308 ( .A(n1157), .B(KEYINPUT72), .ZN(n1160) );
  NAND2_X1 U1309 ( .A1(n1023), .A2(G283), .ZN(n1158) );
  AND2_X1 U1310 ( .A1(n1160), .A2(n1159), .ZN(n1163) );
  NAND2_X1 U1311 ( .A1(G97), .A2(n1466), .ZN(n1161) );
  XOR2_X1 U1312 ( .A(KEYINPUT73), .B(n1161), .Z(n1162) );
  NOR2_X1 U1313 ( .A1(n1214), .A2(n1211), .ZN(n1165) );
  NOR2_X1 U1314 ( .A1(n2043), .A2(n1219), .ZN(n2019) );
  NAND2_X1 U1315 ( .A1(G97), .A2(n1239), .ZN(n1167) );
  NAND2_X1 U1316 ( .A1(G77), .A2(n1466), .ZN(n1166) );
  NAND2_X1 U1317 ( .A1(n1167), .A2(n1166), .ZN(n1172) );
  AND2_X1 U1318 ( .A1(G107), .A2(n1023), .ZN(n1169) );
  NOR2_X1 U1319 ( .A1(G97), .A2(n1462), .ZN(n1168) );
  NOR2_X1 U1320 ( .A1(n1169), .A2(n1168), .ZN(n1170) );
  XNOR2_X1 U1321 ( .A(n1170), .B(KEYINPUT13), .ZN(n1171) );
  NOR2_X1 U1322 ( .A1(n1172), .A2(n1171), .ZN(n1174) );
  XNOR2_X1 U1323 ( .A(G107), .B(G97), .ZN(n2034) );
  NAND2_X1 U1324 ( .A1(n1393), .A2(n2034), .ZN(n1173) );
  NAND2_X1 U1325 ( .A1(n1174), .A2(n1173), .ZN(n1205) );
  AND2_X1 U1326 ( .A1(n1205), .A2(n2043), .ZN(n1175) );
  XOR2_X1 U1327 ( .A(KEYINPUT75), .B(n1175), .Z(n1294) );
  INV_X1 U1328 ( .A(n1188), .ZN(n1187) );
  AND2_X1 U1329 ( .A1(n1180), .A2(n2043), .ZN(n1184) );
  INV_X1 U1330 ( .A(n1211), .ZN(n1182) );
  NAND2_X1 U1331 ( .A1(G200), .A2(n1176), .ZN(n1178) );
  NAND2_X1 U1332 ( .A1(n1178), .A2(n1177), .ZN(n1179) );
  INV_X1 U1333 ( .A(G330), .ZN(n1549) );
  NOR2_X1 U1334 ( .A1(n1796), .A2(n1137), .ZN(n1213) );
  OR2_X1 U1335 ( .A1(n1214), .A2(n1213), .ZN(n1185) );
  NAND2_X1 U1336 ( .A1(n1186), .A2(n1185), .ZN(n1623) );
  NAND2_X1 U1337 ( .A1(n1216), .A2(n1623), .ZN(n2021) );
  NAND2_X1 U1338 ( .A1(n1187), .A2(n2021), .ZN(n1191) );
  INV_X1 U1339 ( .A(n2021), .ZN(n1189) );
  NAND2_X1 U1340 ( .A1(n1189), .A2(n1188), .ZN(n1190) );
  NAND2_X1 U1341 ( .A1(n1191), .A2(n1190), .ZN(n1210) );
  NAND2_X1 U1342 ( .A1(n1434), .A2(G244), .ZN(n1193) );
  NAND2_X1 U1343 ( .A1(n1193), .A2(n1192), .ZN(n1197) );
  NAND2_X1 U1344 ( .A1(G283), .A2(n1444), .ZN(n1195) );
  NAND2_X1 U1345 ( .A1(n1448), .A2(G250), .ZN(n1194) );
  NAND2_X1 U1346 ( .A1(n1195), .A2(n1194), .ZN(n1196) );
  XNOR2_X1 U1347 ( .A(n1199), .B(n1198), .ZN(n1202) );
  NAND2_X1 U1348 ( .A1(n1200), .A2(G257), .ZN(n1201) );
  NAND2_X1 U1349 ( .A1(G200), .A2(n1260), .ZN(n1203) );
  NAND2_X1 U1350 ( .A1(n1203), .A2(n1030), .ZN(n1204) );
  NOR2_X1 U1351 ( .A1(n1205), .A2(n1204), .ZN(n1209) );
  NAND2_X1 U1352 ( .A1(n1441), .A2(n1260), .ZN(n1206) );
  NAND2_X1 U1353 ( .A1(n1206), .A2(n1205), .ZN(n1208) );
  NOR2_X1 U1354 ( .A1(G179), .A2(n1260), .ZN(n1207) );
  NOR2_X1 U1355 ( .A1(n1208), .A2(n1207), .ZN(n1246) );
  NOR2_X1 U1356 ( .A1(n1211), .A2(n2043), .ZN(n1212) );
  NOR2_X1 U1357 ( .A1(n1213), .A2(n1212), .ZN(n1215) );
  XNOR2_X1 U1358 ( .A(n1215), .B(n1214), .ZN(n1217) );
  XNOR2_X1 U1359 ( .A(n1217), .B(n1216), .ZN(n1669) );
  XNOR2_X1 U1360 ( .A(n1218), .B(KEYINPUT52), .ZN(n1782) );
  NAND2_X1 U1361 ( .A1(n1445), .A2(G238), .ZN(n1221) );
  NAND2_X1 U1362 ( .A1(n1448), .A2(G244), .ZN(n1220) );
  NAND2_X1 U1363 ( .A1(n1221), .A2(n1220), .ZN(n1222) );
  XNOR2_X1 U1364 ( .A(n1222), .B(KEYINPUT8), .ZN(n1231) );
  AND2_X1 U1365 ( .A1(G116), .A2(n1444), .ZN(n1226) );
  INV_X1 U1366 ( .A(n1227), .ZN(n1223) );
  NAND2_X1 U1367 ( .A1(G274), .A2(n1223), .ZN(n1224) );
  XOR2_X1 U1368 ( .A(KEYINPUT76), .B(n1224), .Z(n1225) );
  NOR2_X1 U1369 ( .A1(n1226), .A2(n1225), .ZN(n1229) );
  NAND2_X1 U1370 ( .A1(G250), .A2(n1227), .ZN(n1228) );
  NAND2_X1 U1371 ( .A1(n1229), .A2(n1098), .ZN(n1230) );
  NAND2_X1 U1372 ( .A1(G169), .A2(n1259), .ZN(n1233) );
  NAND2_X1 U1373 ( .A1(n1234), .A2(n1233), .ZN(n1795) );
  NOR2_X1 U1374 ( .A1(G87), .A2(n1462), .ZN(n1238) );
  NAND2_X1 U1375 ( .A1(G97), .A2(n1023), .ZN(n1236) );
  NAND2_X1 U1376 ( .A1(G68), .A2(n1466), .ZN(n1235) );
  NAND2_X1 U1377 ( .A1(n1236), .A2(n1235), .ZN(n1237) );
  NOR2_X1 U1378 ( .A1(n1238), .A2(n1237), .ZN(n1245) );
  NOR2_X1 U1379 ( .A1(G107), .A2(G97), .ZN(n1720) );
  INV_X1 U1380 ( .A(G87), .ZN(n1721) );
  NAND2_X1 U1381 ( .A1(n1720), .A2(n1721), .ZN(n1627) );
  NAND2_X1 U1382 ( .A1(G87), .A2(n1239), .ZN(n1241) );
  INV_X1 U1383 ( .A(KEYINPUT78), .ZN(n1240) );
  XNOR2_X1 U1384 ( .A(n1393), .B(n1240), .ZN(n1365) );
  NAND2_X1 U1385 ( .A1(n1241), .A2(n1365), .ZN(n1242) );
  NAND2_X1 U1386 ( .A1(n1627), .A2(n1242), .ZN(n1243) );
  XOR2_X1 U1387 ( .A(KEYINPUT9), .B(n1243), .Z(n1244) );
  NAND2_X1 U1388 ( .A1(n1245), .A2(n1244), .ZN(n1798) );
  INV_X1 U1389 ( .A(n1246), .ZN(n1787) );
  AND2_X1 U1390 ( .A1(n1251), .A2(n1787), .ZN(n1247) );
  INV_X1 U1391 ( .A(n1251), .ZN(n1253) );
  AND2_X1 U1392 ( .A1(n1259), .A2(G200), .ZN(n1248) );
  NOR2_X1 U1393 ( .A1(n1798), .A2(n1248), .ZN(n1250) );
  INV_X1 U1394 ( .A(n1259), .ZN(n1254) );
  NAND2_X1 U1395 ( .A1(G190), .A2(n1254), .ZN(n1249) );
  NAND2_X1 U1396 ( .A1(n1250), .A2(n1249), .ZN(n1790) );
  NAND2_X1 U1397 ( .A1(n1251), .A2(n1790), .ZN(n1252) );
  INV_X1 U1398 ( .A(n1264), .ZN(n1258) );
  NAND2_X1 U1399 ( .A1(n1260), .A2(n1255), .ZN(n1256) );
  NOR2_X1 U1400 ( .A1(n1254), .A2(n1256), .ZN(n1257) );
  NOR2_X1 U1401 ( .A1(n1263), .A2(n1262), .ZN(n1265) );
  AND2_X1 U1402 ( .A1(n1534), .A2(G330), .ZN(n1269) );
  NOR2_X1 U1403 ( .A1(n1293), .A2(n1266), .ZN(n1267) );
  INV_X1 U1404 ( .A(n1283), .ZN(n1275) );
  INV_X1 U1405 ( .A(n1669), .ZN(n1607) );
  NAND2_X1 U1406 ( .A1(n1275), .A2(n1607), .ZN(n1271) );
  NAND2_X1 U1407 ( .A1(n1271), .A2(KEYINPUT79), .ZN(n1272) );
  NOR2_X1 U1408 ( .A1(n2026), .A2(n1272), .ZN(n1273) );
  NOR2_X1 U1409 ( .A1(n1782), .A2(n1273), .ZN(n1278) );
  NOR2_X1 U1410 ( .A1(n1607), .A2(n2026), .ZN(n1274) );
  NOR2_X1 U1411 ( .A1(KEYINPUT79), .A2(n1274), .ZN(n1276) );
  NAND2_X1 U1412 ( .A1(n1276), .A2(n1275), .ZN(n1277) );
  NAND2_X1 U1413 ( .A1(n1287), .A2(n1101), .ZN(n1992) );
  INV_X1 U1414 ( .A(n2031), .ZN(n2023) );
  NAND2_X1 U1415 ( .A1(G45), .A2(n1279), .ZN(n1280) );
  NAND2_X1 U1416 ( .A1(n2022), .A2(n1280), .ZN(n1281) );
  XOR2_X1 U1417 ( .A(KEYINPUT1), .B(n1281), .Z(n1973) );
  INV_X1 U1418 ( .A(n1973), .ZN(n1346) );
  NAND2_X1 U1419 ( .A1(n2031), .A2(n2026), .ZN(n1282) );
  NAND2_X1 U1420 ( .A1(n1346), .A2(n1282), .ZN(n1670) );
  AND2_X1 U1421 ( .A1(n1283), .A2(n1670), .ZN(n1353) );
  INV_X1 U1422 ( .A(n1992), .ZN(n1741) );
  NAND2_X1 U1423 ( .A1(G33), .A2(n1741), .ZN(n1284) );
  XNOR2_X1 U1424 ( .A(n1284), .B(KEYINPUT24), .ZN(n1826) );
  XNOR2_X1 U1425 ( .A(n2034), .B(KEYINPUT51), .ZN(n1286) );
  XNOR2_X1 U1426 ( .A(G87), .B(G116), .ZN(n1285) );
  XNOR2_X1 U1427 ( .A(n1286), .B(n1285), .ZN(n2069) );
  NOR2_X1 U1428 ( .A1(n1826), .A2(n2069), .ZN(n1292) );
  NAND2_X1 U1429 ( .A1(n1287), .A2(n1898), .ZN(n1969) );
  NOR2_X1 U1430 ( .A1(G20), .A2(n1969), .ZN(n1739) );
  NOR2_X1 U1431 ( .A1(G169), .A2(n1121), .ZN(n1288) );
  NOR2_X1 U1432 ( .A1(n1289), .A2(n1288), .ZN(n1572) );
  NOR2_X1 U1433 ( .A1(n1739), .A2(n1572), .ZN(n1823) );
  NAND2_X1 U1434 ( .A1(G97), .A2(n1992), .ZN(n1290) );
  NAND2_X1 U1435 ( .A1(n1823), .A2(n1290), .ZN(n1291) );
  NOR2_X1 U1436 ( .A1(n1292), .A2(n1291), .ZN(n1351) );
  NOR2_X1 U1437 ( .A1(n1294), .A2(n1293), .ZN(n1296) );
  NOR2_X1 U1438 ( .A1(n1787), .A2(n1796), .ZN(n1295) );
  NOR2_X1 U1439 ( .A1(n1296), .A2(n1295), .ZN(n1783) );
  NAND2_X1 U1440 ( .A1(n1783), .A2(n1739), .ZN(n1349) );
  INV_X1 U1441 ( .A(n1572), .ZN(n1883) );
  INV_X1 U1442 ( .A(G200), .ZN(n1417) );
  NAND2_X1 U1443 ( .A1(G190), .A2(n1417), .ZN(n1311) );
  NAND2_X1 U1444 ( .A1(G20), .A2(G179), .ZN(n1297) );
  NAND2_X1 U1445 ( .A1(n1956), .A2(G311), .ZN(n1298) );
  NAND2_X1 U1446 ( .A1(n1298), .A2(G33), .ZN(n1299) );
  XNOR2_X1 U1447 ( .A(n1299), .B(KEYINPUT82), .ZN(n1310) );
  NOR2_X1 U1448 ( .A1(G190), .A2(n1121), .ZN(n1301) );
  NAND2_X1 U1449 ( .A1(G200), .A2(n1301), .ZN(n1302) );
  NAND2_X1 U1450 ( .A1(n1952), .A2(G303), .ZN(n1300) );
  XNOR2_X1 U1451 ( .A(n1300), .B(KEYINPUT84), .ZN(n1308) );
  NAND2_X1 U1452 ( .A1(n1301), .A2(n1417), .ZN(n1303) );
  AND2_X1 U1453 ( .A1(G294), .A2(n1953), .ZN(n1306) );
  NOR2_X1 U1454 ( .A1(G179), .A2(n1302), .ZN(n1832) );
  NAND2_X1 U1455 ( .A1(G107), .A2(n1832), .ZN(n1756) );
  NAND2_X1 U1456 ( .A1(n1943), .A2(G322), .ZN(n1304) );
  NAND2_X1 U1457 ( .A1(n1756), .A2(n1304), .ZN(n1305) );
  NOR2_X1 U1458 ( .A1(n1306), .A2(n1305), .ZN(n1307) );
  NAND2_X1 U1459 ( .A1(n1308), .A2(n1307), .ZN(n1309) );
  NOR2_X1 U1460 ( .A1(n1310), .A2(n1309), .ZN(n1315) );
  OR2_X1 U1461 ( .A1(n1311), .A2(G179), .ZN(n1312) );
  NAND2_X1 U1462 ( .A1(n1312), .A2(G20), .ZN(n1313) );
  XOR2_X1 U1463 ( .A(KEYINPUT83), .B(n1313), .Z(n1860) );
  NAND2_X1 U1464 ( .A1(G116), .A2(n1860), .ZN(n1314) );
  NAND2_X1 U1465 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
  XNOR2_X1 U1466 ( .A(KEYINPUT58), .B(n1316), .ZN(n1325) );
  NAND2_X1 U1467 ( .A1(G200), .A2(G190), .ZN(n1317) );
  XOR2_X1 U1468 ( .A(KEYINPUT80), .B(n1317), .Z(n1318) );
  NAND2_X1 U1469 ( .A1(G20), .A2(n1318), .ZN(n1319) );
  NAND2_X1 U1470 ( .A1(G317), .A2(n1947), .ZN(n1321) );
  NAND2_X1 U1471 ( .A1(n1946), .A2(G283), .ZN(n1320) );
  NAND2_X1 U1472 ( .A1(n1321), .A2(n1320), .ZN(n1322) );
  XNOR2_X1 U1473 ( .A(KEYINPUT81), .B(n1322), .ZN(n1323) );
  XNOR2_X1 U1474 ( .A(KEYINPUT59), .B(n1323), .ZN(n1324) );
  NOR2_X1 U1475 ( .A1(n1325), .A2(n1324), .ZN(n1344) );
  INV_X1 U1476 ( .A(n1860), .ZN(n1932) );
  INV_X1 U1477 ( .A(G77), .ZN(n2054) );
  NOR2_X1 U1478 ( .A1(n1932), .A2(n2054), .ZN(n1703) );
  NAND2_X1 U1479 ( .A1(n1832), .A2(G87), .ZN(n1326) );
  XNOR2_X1 U1480 ( .A(n1326), .B(KEYINPUT22), .ZN(n1885) );
  NAND2_X1 U1481 ( .A1(n1956), .A2(G159), .ZN(n1327) );
  NAND2_X1 U1482 ( .A1(n1898), .A2(n1327), .ZN(n1331) );
  NAND2_X1 U1483 ( .A1(G50), .A2(n1952), .ZN(n1329) );
  NAND2_X1 U1484 ( .A1(G143), .A2(n1943), .ZN(n1328) );
  NAND2_X1 U1485 ( .A1(n1329), .A2(n1328), .ZN(n1330) );
  NOR2_X1 U1486 ( .A1(n1331), .A2(n1330), .ZN(n1333) );
  NAND2_X1 U1487 ( .A1(n1953), .A2(G58), .ZN(n1332) );
  NAND2_X1 U1488 ( .A1(n1333), .A2(n1332), .ZN(n1340) );
  NAND2_X1 U1489 ( .A1(n1947), .A2(G150), .ZN(n1334) );
  XNOR2_X1 U1490 ( .A(n1334), .B(KEYINPUT56), .ZN(n1336) );
  NAND2_X1 U1491 ( .A1(n1946), .A2(G68), .ZN(n1335) );
  NAND2_X1 U1492 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
  XNOR2_X1 U1493 ( .A(KEYINPUT85), .B(n1337), .ZN(n1338) );
  XNOR2_X1 U1494 ( .A(KEYINPUT57), .B(n1338), .ZN(n1339) );
  NOR2_X1 U1495 ( .A1(n1340), .A2(n1339), .ZN(n1341) );
  NAND2_X1 U1496 ( .A1(n1885), .A2(n1341), .ZN(n1342) );
  NOR2_X1 U1497 ( .A1(n1703), .A2(n1342), .ZN(n1343) );
  NOR2_X1 U1498 ( .A1(n1344), .A2(n1343), .ZN(n1345) );
  NOR2_X1 U1499 ( .A1(n1883), .A2(n1345), .ZN(n1347) );
  NAND2_X1 U1500 ( .A1(n1346), .A2(n2023), .ZN(n1940) );
  NOR2_X1 U1501 ( .A1(n1347), .A2(n1940), .ZN(n1348) );
  NAND2_X1 U1502 ( .A1(n1349), .A2(n1348), .ZN(n1350) );
  NOR2_X1 U1503 ( .A1(n1351), .A2(n1350), .ZN(n1352) );
  OR2_X1 U1504 ( .A1(n1353), .A2(n1352), .ZN(n1354) );
  NAND2_X1 U1505 ( .A1(n1023), .A2(G58), .ZN(n1358) );
  INV_X1 U1506 ( .A(G50), .ZN(n2063) );
  NAND2_X1 U1507 ( .A1(n1356), .A2(n2063), .ZN(n1357) );
  NAND2_X1 U1508 ( .A1(n1358), .A2(n1357), .ZN(n1362) );
  NOR2_X1 U1509 ( .A1(n1360), .A2(n1359), .ZN(n1423) );
  NOR2_X1 U1510 ( .A1(n1423), .A2(n1393), .ZN(n1469) );
  NOR2_X1 U1511 ( .A1(n1469), .A2(n2063), .ZN(n1361) );
  NOR2_X1 U1512 ( .A1(n1362), .A2(n1361), .ZN(n1364) );
  NAND2_X1 U1513 ( .A1(n1466), .A2(G150), .ZN(n1363) );
  NAND2_X1 U1514 ( .A1(n1364), .A2(n1363), .ZN(n1367) );
  NOR2_X1 U1515 ( .A1(G68), .A2(G58), .ZN(n2064) );
  NOR2_X1 U1516 ( .A1(n2064), .A2(n1365), .ZN(n1366) );
  NOR2_X1 U1517 ( .A1(n1367), .A2(n1366), .ZN(n1552) );
  NAND2_X1 U1518 ( .A1(n1448), .A2(G223), .ZN(n1369) );
  NAND2_X1 U1519 ( .A1(G77), .A2(n1444), .ZN(n1368) );
  NAND2_X1 U1520 ( .A1(n1369), .A2(n1368), .ZN(n1375) );
  NOR2_X1 U1521 ( .A1(G45), .A2(G41), .ZN(n1370) );
  NOR2_X1 U1522 ( .A1(n2022), .A2(n1370), .ZN(n1371) );
  NAND2_X1 U1523 ( .A1(G274), .A2(n1371), .ZN(n1453) );
  NOR2_X1 U1524 ( .A1(n1372), .A2(n1371), .ZN(n1456) );
  NAND2_X1 U1525 ( .A1(n1456), .A2(G226), .ZN(n1373) );
  NAND2_X1 U1526 ( .A1(n1453), .A2(n1373), .ZN(n1374) );
  XOR2_X1 U1527 ( .A(KEYINPUT98), .B(n1376), .Z(n1380) );
  NAND2_X1 U1528 ( .A1(G222), .A2(n1434), .ZN(n1378) );
  NAND2_X1 U1529 ( .A1(G190), .A2(n1386), .ZN(n1383) );
  NAND2_X1 U1530 ( .A1(n1552), .A2(n1383), .ZN(n1385) );
  NOR2_X1 U1531 ( .A1(n1386), .A2(n1417), .ZN(n1384) );
  NOR2_X1 U1532 ( .A1(n1385), .A2(n1384), .ZN(n1389) );
  NOR2_X1 U1533 ( .A1(n1027), .A2(n1552), .ZN(n1388) );
  OR2_X1 U1534 ( .A1(G169), .A2(n1386), .ZN(n1387) );
  XNOR2_X1 U1535 ( .A(n1390), .B(KEYINPUT37), .ZN(n1483) );
  NAND2_X1 U1536 ( .A1(G159), .A2(n1466), .ZN(n1399) );
  NAND2_X1 U1537 ( .A1(n1023), .A2(G68), .ZN(n1392) );
  OR2_X1 U1538 ( .A1(n1462), .A2(G58), .ZN(n1391) );
  NAND2_X1 U1539 ( .A1(n1392), .A2(n1391), .ZN(n1397) );
  NAND2_X1 U1540 ( .A1(n1423), .A2(G58), .ZN(n1395) );
  XNOR2_X1 U1541 ( .A(G68), .B(G58), .ZN(n1743) );
  NAND2_X1 U1542 ( .A1(n1743), .A2(n1393), .ZN(n1394) );
  NAND2_X1 U1543 ( .A1(n1395), .A2(n1394), .ZN(n1396) );
  NOR2_X1 U1544 ( .A1(n1397), .A2(n1396), .ZN(n1398) );
  NAND2_X1 U1545 ( .A1(n1399), .A2(n1398), .ZN(n1400) );
  XNOR2_X1 U1546 ( .A(n1400), .B(KEYINPUT30), .ZN(n1521) );
  NAND2_X1 U1547 ( .A1(n1444), .A2(G87), .ZN(n1401) );
  XOR2_X1 U1548 ( .A(KEYINPUT31), .B(n1401), .Z(n1403) );
  NAND2_X1 U1549 ( .A1(n1456), .A2(G232), .ZN(n1402) );
  NAND2_X1 U1550 ( .A1(n1403), .A2(n1402), .ZN(n1410) );
  NAND2_X1 U1551 ( .A1(n1448), .A2(G226), .ZN(n1404) );
  XNOR2_X1 U1552 ( .A(n1404), .B(KEYINPUT32), .ZN(n1406) );
  NAND2_X1 U1553 ( .A1(G223), .A2(n1434), .ZN(n1405) );
  NAND2_X1 U1554 ( .A1(n1406), .A2(n1405), .ZN(n1407) );
  XNOR2_X1 U1555 ( .A(n1407), .B(KEYINPUT33), .ZN(n1408) );
  NAND2_X1 U1556 ( .A1(n1408), .A2(n1453), .ZN(n1409) );
  NOR2_X2 U1557 ( .A1(n1410), .A2(n1409), .ZN(n1419) );
  INV_X1 U1558 ( .A(n1419), .ZN(n1413) );
  XNOR2_X1 U1559 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n1411) );
  XNOR2_X1 U1560 ( .A(n1412), .B(n1411), .ZN(n1415) );
  NAND2_X1 U1561 ( .A1(n1413), .A2(G169), .ZN(n1414) );
  NAND2_X1 U1562 ( .A1(n1415), .A2(n1414), .ZN(n1416) );
  NOR2_X1 U1563 ( .A1(n1419), .A2(n1417), .ZN(n1418) );
  XNOR2_X1 U1564 ( .A(n1418), .B(KEYINPUT35), .ZN(n1421) );
  NAND2_X1 U1565 ( .A1(n1419), .A2(G190), .ZN(n1420) );
  NAND2_X1 U1566 ( .A1(n1421), .A2(n1420), .ZN(n1422) );
  NOR2_X1 U1567 ( .A1(n1521), .A2(n1422), .ZN(n1484) );
  NAND2_X1 U1568 ( .A1(n1423), .A2(G68), .ZN(n1424) );
  XNOR2_X1 U1569 ( .A(n1424), .B(KEYINPUT93), .ZN(n1426) );
  INV_X1 U1570 ( .A(n1023), .ZN(n1463) );
  NOR2_X1 U1571 ( .A1(n2054), .A2(n1463), .ZN(n1425) );
  NOR2_X1 U1572 ( .A1(n1426), .A2(n1425), .ZN(n1428) );
  NAND2_X1 U1573 ( .A1(n1466), .A2(G50), .ZN(n1427) );
  NAND2_X1 U1574 ( .A1(n1428), .A2(n1427), .ZN(n1431) );
  NOR2_X1 U1575 ( .A1(n1429), .A2(G68), .ZN(n1430) );
  NAND2_X1 U1576 ( .A1(n1456), .A2(G238), .ZN(n1432) );
  XNOR2_X1 U1577 ( .A(n1432), .B(KEYINPUT94), .ZN(n1440) );
  NAND2_X1 U1578 ( .A1(G97), .A2(n1444), .ZN(n1433) );
  NAND2_X1 U1579 ( .A1(n1453), .A2(n1433), .ZN(n1438) );
  NAND2_X1 U1580 ( .A1(n1434), .A2(G226), .ZN(n1436) );
  NAND2_X1 U1581 ( .A1(n1448), .A2(G232), .ZN(n1435) );
  NAND2_X1 U1582 ( .A1(n1436), .A2(n1435), .ZN(n1437) );
  XNOR2_X1 U1583 ( .A(n1017), .B(KEYINPUT95), .ZN(n1443) );
  NAND2_X1 U1584 ( .A1(G107), .A2(n1444), .ZN(n1447) );
  NAND2_X1 U1585 ( .A1(G232), .A2(n1445), .ZN(n1446) );
  NAND2_X1 U1586 ( .A1(n1447), .A2(n1446), .ZN(n1452) );
  NAND2_X1 U1587 ( .A1(n1448), .A2(G238), .ZN(n1450) );
  XNOR2_X1 U1588 ( .A(n1450), .B(n1449), .ZN(n1451) );
  NOR2_X1 U1589 ( .A1(n1452), .A2(n1451), .ZN(n1454) );
  NAND2_X1 U1590 ( .A1(n1454), .A2(n1453), .ZN(n1455) );
  XNOR2_X1 U1591 ( .A(n1455), .B(KEYINPUT7), .ZN(n1458) );
  NAND2_X1 U1592 ( .A1(n1456), .A2(G244), .ZN(n1457) );
  NAND2_X1 U1593 ( .A1(n1458), .A2(n1457), .ZN(n1485) );
  NOR2_X1 U1594 ( .A1(n1084), .A2(n1485), .ZN(n1460) );
  AND2_X1 U1595 ( .A1(n1485), .A2(G169), .ZN(n1459) );
  NOR2_X1 U1596 ( .A1(n1460), .A2(n1459), .ZN(n1461) );
  XNOR2_X1 U1597 ( .A(n1461), .B(KEYINPUT92), .ZN(n1512) );
  NOR2_X1 U1598 ( .A1(G77), .A2(n1462), .ZN(n1465) );
  NOR2_X1 U1599 ( .A1(n1463), .A2(n1721), .ZN(n1464) );
  NOR2_X1 U1600 ( .A1(n1465), .A2(n1464), .ZN(n1468) );
  NAND2_X1 U1601 ( .A1(n1466), .A2(G58), .ZN(n1467) );
  NAND2_X1 U1602 ( .A1(n1468), .A2(n1467), .ZN(n1471) );
  NOR2_X1 U1603 ( .A1(n1469), .A2(n2054), .ZN(n1470) );
  NOR2_X1 U1604 ( .A1(n1471), .A2(n1470), .ZN(n1508) );
  XOR2_X1 U1605 ( .A(KEYINPUT28), .B(n1472), .Z(n1476) );
  XNOR2_X1 U1606 ( .A(n1473), .B(KEYINPUT27), .ZN(n1474) );
  NOR2_X1 U1607 ( .A1(n1474), .A2(n1015), .ZN(n1475) );
  NAND2_X1 U1608 ( .A1(n1476), .A2(n1475), .ZN(n1477) );
  NOR2_X1 U1609 ( .A1(n1498), .A2(n1500), .ZN(n1478) );
  NOR2_X1 U1610 ( .A1(n1501), .A2(n1478), .ZN(n1479) );
  NOR2_X1 U1611 ( .A1(n1484), .A2(n1479), .ZN(n1480) );
  NOR2_X1 U1612 ( .A1(n1542), .A2(n1480), .ZN(n1481) );
  NOR2_X1 U1613 ( .A1(n1483), .A2(n1481), .ZN(n1482) );
  NOR2_X1 U1614 ( .A1(n1500), .A2(n1483), .ZN(n1492) );
  XNOR2_X1 U1615 ( .A(KEYINPUT91), .B(n1508), .ZN(n1487) );
  NOR2_X1 U1616 ( .A1(n1083), .A2(n1485), .ZN(n1486) );
  NOR2_X1 U1617 ( .A1(n1487), .A2(n1486), .ZN(n1489) );
  NAND2_X1 U1618 ( .A1(G200), .A2(n1485), .ZN(n1488) );
  NAND2_X1 U1619 ( .A1(n1489), .A2(n1488), .ZN(n1496) );
  NAND2_X1 U1620 ( .A1(n2042), .A2(n1493), .ZN(G369) );
  NOR2_X1 U1621 ( .A1(n2043), .A2(n1494), .ZN(n1507) );
  OR2_X1 U1622 ( .A1(n2043), .A2(n1498), .ZN(n1499) );
  NAND2_X1 U1623 ( .A1(n1501), .A2(n2043), .ZN(n1502) );
  XOR2_X1 U1624 ( .A(KEYINPUT96), .B(KEYINPUT29), .Z(n1504) );
  NOR2_X1 U1625 ( .A1(n1529), .A2(n1531), .ZN(n1506) );
  NOR2_X1 U1626 ( .A1(n1508), .A2(n1796), .ZN(n1509) );
  XOR2_X1 U1627 ( .A(KEYINPUT5), .B(n1509), .Z(n1511) );
  NOR2_X1 U1628 ( .A1(n1511), .A2(n1510), .ZN(n1515) );
  INV_X1 U1629 ( .A(n1511), .ZN(n1513) );
  NOR2_X1 U1630 ( .A1(n1513), .A2(n1512), .ZN(n1514) );
  NOR2_X1 U1631 ( .A1(n1515), .A2(n1514), .ZN(n1903) );
  INV_X1 U1632 ( .A(n1903), .ZN(n1517) );
  INV_X1 U1633 ( .A(n1531), .ZN(n1516) );
  NAND2_X1 U1634 ( .A1(n1517), .A2(n1516), .ZN(n1518) );
  XNOR2_X1 U1635 ( .A(n1519), .B(KEYINPUT39), .ZN(n1520) );
  NAND2_X1 U1636 ( .A1(n1521), .A2(n1555), .ZN(n1523) );
  NAND2_X1 U1637 ( .A1(n1523), .A2(n1522), .ZN(n1525) );
  NAND2_X1 U1638 ( .A1(n1542), .A2(n1555), .ZN(n1524) );
  NAND2_X1 U1639 ( .A1(n1530), .A2(n1529), .ZN(n1532) );
  XNOR2_X2 U1640 ( .A(n1532), .B(n1531), .ZN(n1972) );
  AND2_X1 U1641 ( .A1(n1534), .A2(n1533), .ZN(n1548) );
  NAND2_X1 U1642 ( .A1(n1548), .A2(n2018), .ZN(n2040) );
  NOR2_X1 U1643 ( .A1(n1549), .A2(n2040), .ZN(n1535) );
  NOR2_X1 U1644 ( .A1(G369), .A2(n1535), .ZN(n1537) );
  XNOR2_X1 U1645 ( .A(n1537), .B(n1536), .ZN(n1919) );
  NOR2_X1 U1646 ( .A1(n1919), .A2(n1973), .ZN(n1538) );
  INV_X1 U1647 ( .A(n1540), .ZN(n1541) );
  NAND2_X1 U1648 ( .A1(n1674), .A2(n1541), .ZN(n1544) );
  INV_X1 U1649 ( .A(n1555), .ZN(n1551) );
  NAND2_X1 U1650 ( .A1(n1542), .A2(n1551), .ZN(n1543) );
  NAND2_X1 U1651 ( .A1(n1544), .A2(n1543), .ZN(n2045) );
  XNOR2_X1 U1652 ( .A(KEYINPUT100), .B(n1674), .ZN(n1545) );
  NAND2_X1 U1653 ( .A1(n1545), .A2(n1516), .ZN(n1546) );
  NOR2_X1 U1654 ( .A1(n1903), .A2(n1546), .ZN(n1547) );
  NAND2_X1 U1655 ( .A1(n1548), .A2(n1547), .ZN(n2039) );
  NOR2_X1 U1656 ( .A1(n1549), .A2(n2039), .ZN(n1550) );
  NOR2_X1 U1657 ( .A1(n2045), .A2(n1550), .ZN(n1559) );
  OR2_X1 U1658 ( .A1(n1552), .A2(n1551), .ZN(n1554) );
  INV_X1 U1659 ( .A(n1483), .ZN(n1553) );
  NAND2_X1 U1660 ( .A1(n1554), .A2(n1553), .ZN(n1558) );
  NAND2_X1 U1661 ( .A1(n1556), .A2(n1555), .ZN(n1557) );
  NAND2_X1 U1662 ( .A1(n1558), .A2(n1557), .ZN(n1563) );
  XNOR2_X1 U1663 ( .A(n1559), .B(n1563), .ZN(n1560) );
  INV_X1 U1664 ( .A(n1940), .ZN(n1859) );
  OR2_X1 U1665 ( .A1(n1883), .A2(G41), .ZN(n1561) );
  NAND2_X1 U1666 ( .A1(n1561), .A2(n2063), .ZN(n1562) );
  NAND2_X1 U1667 ( .A1(n1969), .A2(n1562), .ZN(n1565) );
  INV_X1 U1668 ( .A(n1969), .ZN(n1902) );
  NAND2_X1 U1669 ( .A1(n1902), .A2(n1563), .ZN(n1564) );
  NAND2_X1 U1670 ( .A1(n1565), .A2(n1564), .ZN(n1604) );
  NAND2_X1 U1671 ( .A1(G87), .A2(n1953), .ZN(n1566) );
  XNOR2_X1 U1672 ( .A(n1566), .B(KEYINPUT102), .ZN(n1567) );
  NAND2_X1 U1673 ( .A1(G68), .A2(n1860), .ZN(n1831) );
  NAND2_X1 U1674 ( .A1(n1567), .A2(n1831), .ZN(n1580) );
  NAND2_X1 U1675 ( .A1(n1832), .A2(G58), .ZN(n1927) );
  NAND2_X1 U1676 ( .A1(G283), .A2(n1943), .ZN(n1568) );
  NAND2_X1 U1677 ( .A1(n1927), .A2(n1568), .ZN(n1571) );
  NAND2_X1 U1678 ( .A1(G107), .A2(n1956), .ZN(n1569) );
  XOR2_X1 U1679 ( .A(KEYINPUT42), .B(n1569), .Z(n1570) );
  NOR2_X1 U1680 ( .A1(n1571), .A2(n1570), .ZN(n1578) );
  INV_X1 U1681 ( .A(n1946), .ZN(n1697) );
  NOR2_X1 U1682 ( .A1(n2054), .A2(n1697), .ZN(n1619) );
  NAND2_X1 U1683 ( .A1(G33), .A2(n1572), .ZN(n1941) );
  NOR2_X1 U1684 ( .A1(n1619), .A2(n1941), .ZN(n1574) );
  NAND2_X1 U1685 ( .A1(G97), .A2(n1952), .ZN(n1573) );
  NAND2_X1 U1686 ( .A1(n1574), .A2(n1573), .ZN(n1576) );
  AND2_X1 U1687 ( .A1(G116), .A2(n1947), .ZN(n1575) );
  NOR2_X1 U1688 ( .A1(n1576), .A2(n1575), .ZN(n1577) );
  NAND2_X1 U1689 ( .A1(n1578), .A2(n1577), .ZN(n1579) );
  NOR2_X1 U1690 ( .A1(n1580), .A2(n1579), .ZN(n1600) );
  NOR2_X1 U1691 ( .A1(G33), .A2(n1883), .ZN(n1931) );
  INV_X1 U1692 ( .A(n1931), .ZN(n1677) );
  NAND2_X1 U1693 ( .A1(G128), .A2(n1956), .ZN(n1582) );
  NAND2_X1 U1694 ( .A1(G124), .A2(n1943), .ZN(n1581) );
  NAND2_X1 U1695 ( .A1(n1582), .A2(n1581), .ZN(n1583) );
  NOR2_X1 U1696 ( .A1(n1677), .A2(n1583), .ZN(n1593) );
  NAND2_X1 U1697 ( .A1(G143), .A2(n1946), .ZN(n1585) );
  NAND2_X1 U1698 ( .A1(G125), .A2(n1947), .ZN(n1584) );
  NAND2_X1 U1699 ( .A1(n1585), .A2(n1584), .ZN(n1591) );
  NAND2_X1 U1700 ( .A1(n1952), .A2(G132), .ZN(n1586) );
  XOR2_X1 U1701 ( .A(KEYINPUT101), .B(n1586), .Z(n1588) );
  NAND2_X1 U1702 ( .A1(n1832), .A2(G159), .ZN(n1587) );
  NAND2_X1 U1703 ( .A1(n1588), .A2(n1587), .ZN(n1589) );
  XNOR2_X1 U1704 ( .A(KEYINPUT44), .B(n1589), .ZN(n1590) );
  NOR2_X1 U1705 ( .A1(n1591), .A2(n1590), .ZN(n1592) );
  NAND2_X1 U1706 ( .A1(n1593), .A2(n1592), .ZN(n1598) );
  NAND2_X1 U1707 ( .A1(G137), .A2(n1953), .ZN(n1594) );
  XOR2_X1 U1708 ( .A(KEYINPUT43), .B(n1594), .Z(n1596) );
  NAND2_X1 U1709 ( .A1(G150), .A2(n1860), .ZN(n1595) );
  NAND2_X1 U1710 ( .A1(n1596), .A2(n1595), .ZN(n1597) );
  NOR2_X1 U1711 ( .A1(n1598), .A2(n1597), .ZN(n1599) );
  NOR2_X1 U1712 ( .A1(n1600), .A2(n1599), .ZN(n1601) );
  NOR2_X1 U1713 ( .A1(G41), .A2(n1601), .ZN(n1602) );
  NOR2_X1 U1714 ( .A1(n1602), .A2(n1940), .ZN(n1603) );
  NAND2_X1 U1715 ( .A1(n1604), .A2(n1603), .ZN(n1605) );
  NOR2_X1 U1716 ( .A1(n2023), .A2(n2026), .ZN(n1606) );
  NAND2_X1 U1717 ( .A1(n1607), .A2(n1606), .ZN(n1608) );
  XNOR2_X1 U1718 ( .A(n1608), .B(KEYINPUT109), .ZN(n1667) );
  NAND2_X1 U1719 ( .A1(G159), .A2(n1947), .ZN(n1621) );
  NAND2_X1 U1720 ( .A1(G50), .A2(n1956), .ZN(n1610) );
  NAND2_X1 U1721 ( .A1(G150), .A2(n1943), .ZN(n1609) );
  NAND2_X1 U1722 ( .A1(n1610), .A2(n1609), .ZN(n1613) );
  NAND2_X1 U1723 ( .A1(G97), .A2(n1832), .ZN(n1804) );
  NAND2_X1 U1724 ( .A1(G68), .A2(n1953), .ZN(n1611) );
  NAND2_X1 U1725 ( .A1(n1804), .A2(n1611), .ZN(n1612) );
  NOR2_X1 U1726 ( .A1(n1613), .A2(n1612), .ZN(n1617) );
  NOR2_X1 U1727 ( .A1(n1932), .A2(n1721), .ZN(n1942) );
  NAND2_X1 U1728 ( .A1(n1952), .A2(G58), .ZN(n1614) );
  NAND2_X1 U1729 ( .A1(n1931), .A2(n1614), .ZN(n1615) );
  NOR2_X1 U1730 ( .A1(n1942), .A2(n1615), .ZN(n1616) );
  NAND2_X1 U1731 ( .A1(n1617), .A2(n1616), .ZN(n1618) );
  NOR2_X1 U1732 ( .A1(n1619), .A2(n1618), .ZN(n1620) );
  NAND2_X1 U1733 ( .A1(n1621), .A2(n1620), .ZN(n1622) );
  NAND2_X1 U1734 ( .A1(n1622), .A2(n1859), .ZN(n1625) );
  INV_X1 U1735 ( .A(n1739), .ZN(n1846) );
  NOR2_X1 U1736 ( .A1(n1623), .A2(n1846), .ZN(n1624) );
  NOR2_X1 U1737 ( .A1(n1625), .A2(n1624), .ZN(n1645) );
  NOR2_X1 U1738 ( .A1(n1741), .A2(G107), .ZN(n1626) );
  XNOR2_X1 U1739 ( .A(KEYINPUT107), .B(n1626), .ZN(n1642) );
  NOR2_X1 U1740 ( .A1(G116), .A2(n1627), .ZN(n2024) );
  NAND2_X1 U1741 ( .A1(G77), .A2(G68), .ZN(n1628) );
  NAND2_X1 U1742 ( .A1(n2024), .A2(n1628), .ZN(n1630) );
  NAND2_X1 U1743 ( .A1(G58), .A2(n2063), .ZN(n1629) );
  NOR2_X1 U1744 ( .A1(n1630), .A2(n1629), .ZN(n1631) );
  NOR2_X1 U1745 ( .A1(G45), .A2(n1631), .ZN(n1632) );
  XOR2_X1 U1746 ( .A(KEYINPUT23), .B(n1632), .Z(n1637) );
  INV_X1 U1747 ( .A(G45), .ZN(n1745) );
  XOR2_X1 U1748 ( .A(KEYINPUT108), .B(G226), .Z(n1634) );
  XNOR2_X1 U1749 ( .A(G244), .B(G238), .ZN(n1633) );
  XNOR2_X1 U1750 ( .A(n1634), .B(n1633), .ZN(n1635) );
  XOR2_X1 U1751 ( .A(G232), .B(n1635), .Z(n2066) );
  NOR2_X1 U1752 ( .A1(n1745), .A2(n2066), .ZN(n1636) );
  NOR2_X1 U1753 ( .A1(n1637), .A2(n1636), .ZN(n1638) );
  NOR2_X1 U1754 ( .A1(n1826), .A2(n1638), .ZN(n1640) );
  NOR2_X1 U1755 ( .A1(n2024), .A2(n1969), .ZN(n1639) );
  NOR2_X1 U1756 ( .A1(n1640), .A2(n1639), .ZN(n1641) );
  NAND2_X1 U1757 ( .A1(n1642), .A2(n1641), .ZN(n1643) );
  NAND2_X1 U1758 ( .A1(n1643), .A2(n1823), .ZN(n1644) );
  NAND2_X1 U1759 ( .A1(n1645), .A2(n1644), .ZN(n1665) );
  NAND2_X1 U1760 ( .A1(G322), .A2(n1947), .ZN(n1647) );
  NAND2_X1 U1761 ( .A1(n1946), .A2(G294), .ZN(n1646) );
  NAND2_X1 U1762 ( .A1(n1647), .A2(n1646), .ZN(n1648) );
  XNOR2_X1 U1763 ( .A(KEYINPUT26), .B(n1648), .ZN(n1663) );
  NAND2_X1 U1764 ( .A1(G326), .A2(n1943), .ZN(n1650) );
  NAND2_X1 U1765 ( .A1(n1952), .A2(G311), .ZN(n1649) );
  NAND2_X1 U1766 ( .A1(n1650), .A2(n1649), .ZN(n1658) );
  NAND2_X1 U1767 ( .A1(n1956), .A2(G317), .ZN(n1652) );
  NAND2_X1 U1768 ( .A1(n1953), .A2(G303), .ZN(n1651) );
  NAND2_X1 U1769 ( .A1(n1652), .A2(n1651), .ZN(n1653) );
  NOR2_X1 U1770 ( .A1(n1941), .A2(n1653), .ZN(n1656) );
  NAND2_X1 U1771 ( .A1(n1832), .A2(G116), .ZN(n1654) );
  XOR2_X1 U1772 ( .A(KEYINPUT25), .B(n1654), .Z(n1655) );
  NAND2_X1 U1773 ( .A1(n1656), .A2(n1655), .ZN(n1657) );
  NOR2_X1 U1774 ( .A1(n1658), .A2(n1657), .ZN(n1660) );
  NAND2_X1 U1775 ( .A1(G283), .A2(n1860), .ZN(n1659) );
  NAND2_X1 U1776 ( .A1(n1660), .A2(n1659), .ZN(n1661) );
  XNOR2_X1 U1777 ( .A(KEYINPUT106), .B(n1661), .ZN(n1662) );
  NOR2_X1 U1778 ( .A1(n1663), .A2(n1662), .ZN(n1664) );
  NOR2_X1 U1779 ( .A1(n1665), .A2(n1664), .ZN(n1666) );
  XNOR2_X1 U1780 ( .A(n1668), .B(KEYINPUT110), .ZN(n1672) );
  NAND2_X1 U1781 ( .A1(n1670), .A2(n1669), .ZN(n1671) );
  NAND2_X1 U1782 ( .A1(n1672), .A2(n1671), .ZN(G393) );
  NAND2_X1 U1783 ( .A1(n1969), .A2(n1883), .ZN(n1965) );
  NOR2_X1 U1784 ( .A1(G58), .A2(n1965), .ZN(n1673) );
  NOR2_X1 U1785 ( .A1(n1940), .A2(n1673), .ZN(n1696) );
  NOR2_X1 U1786 ( .A1(n1969), .A2(n1674), .ZN(n1694) );
  NAND2_X1 U1787 ( .A1(n1946), .A2(G150), .ZN(n1675) );
  XNOR2_X1 U1788 ( .A(KEYINPUT103), .B(n1675), .ZN(n1676) );
  NOR2_X1 U1789 ( .A1(n1677), .A2(n1676), .ZN(n1678) );
  XNOR2_X1 U1790 ( .A(n1678), .B(KEYINPUT104), .ZN(n1680) );
  NAND2_X1 U1791 ( .A1(G128), .A2(n1947), .ZN(n1679) );
  NAND2_X1 U1792 ( .A1(n1680), .A2(n1679), .ZN(n1692) );
  NAND2_X1 U1793 ( .A1(G137), .A2(n1952), .ZN(n1682) );
  NAND2_X1 U1794 ( .A1(G125), .A2(n1943), .ZN(n1681) );
  NAND2_X1 U1795 ( .A1(n1682), .A2(n1681), .ZN(n1684) );
  AND2_X1 U1796 ( .A1(n1860), .A2(G159), .ZN(n1683) );
  NOR2_X1 U1797 ( .A1(n1684), .A2(n1683), .ZN(n1690) );
  NAND2_X1 U1798 ( .A1(G132), .A2(n1956), .ZN(n1686) );
  NAND2_X1 U1799 ( .A1(G143), .A2(n1953), .ZN(n1685) );
  NAND2_X1 U1800 ( .A1(n1686), .A2(n1685), .ZN(n1688) );
  AND2_X1 U1801 ( .A1(n1832), .A2(G50), .ZN(n1687) );
  NOR2_X1 U1802 ( .A1(n1688), .A2(n1687), .ZN(n1689) );
  NAND2_X1 U1803 ( .A1(n1690), .A2(n1689), .ZN(n1691) );
  NOR2_X1 U1804 ( .A1(n1692), .A2(n1691), .ZN(n1693) );
  NOR2_X1 U1805 ( .A1(n1694), .A2(n1693), .ZN(n1695) );
  NAND2_X1 U1806 ( .A1(n1696), .A2(n1695), .ZN(n1714) );
  NOR2_X1 U1807 ( .A1(n1721), .A2(n1697), .ZN(n1773) );
  NAND2_X1 U1808 ( .A1(n1953), .A2(G97), .ZN(n1699) );
  NAND2_X1 U1809 ( .A1(n1943), .A2(G294), .ZN(n1698) );
  NAND2_X1 U1810 ( .A1(n1699), .A2(n1698), .ZN(n1700) );
  XNOR2_X1 U1811 ( .A(KEYINPUT48), .B(n1700), .ZN(n1707) );
  NAND2_X1 U1812 ( .A1(G68), .A2(n1832), .ZN(n1875) );
  NAND2_X1 U1813 ( .A1(G107), .A2(n1952), .ZN(n1701) );
  NAND2_X1 U1814 ( .A1(n1875), .A2(n1701), .ZN(n1702) );
  NOR2_X1 U1815 ( .A1(n1703), .A2(n1702), .ZN(n1705) );
  NAND2_X1 U1816 ( .A1(G283), .A2(n1947), .ZN(n1704) );
  NAND2_X1 U1817 ( .A1(n1705), .A2(n1704), .ZN(n1706) );
  NOR2_X1 U1818 ( .A1(n1707), .A2(n1706), .ZN(n1711) );
  NAND2_X1 U1819 ( .A1(n1956), .A2(G116), .ZN(n1708) );
  XNOR2_X1 U1820 ( .A(KEYINPUT47), .B(n1708), .ZN(n1709) );
  NOR2_X1 U1821 ( .A1(n1941), .A2(n1709), .ZN(n1710) );
  NAND2_X1 U1822 ( .A1(n1711), .A2(n1710), .ZN(n1712) );
  NOR2_X1 U1823 ( .A1(n1773), .A2(n1712), .ZN(n1713) );
  INV_X1 U1824 ( .A(n1919), .ZN(n1716) );
  NAND2_X1 U1825 ( .A1(n1716), .A2(n1972), .ZN(n1717) );
  XNOR2_X1 U1826 ( .A(n1715), .B(n1717), .ZN(n1718) );
  NAND2_X1 U1827 ( .A1(n1715), .A2(n1973), .ZN(n1719) );
  OR2_X1 U1828 ( .A1(n1721), .A2(n1720), .ZN(G355) );
  XNOR2_X1 U1829 ( .A(n1022), .B(G330), .ZN(n1722) );
  NAND2_X1 U1830 ( .A1(n1722), .A2(n1940), .ZN(n1781) );
  NAND2_X1 U1831 ( .A1(G303), .A2(n1946), .ZN(n1738) );
  NAND2_X1 U1832 ( .A1(G283), .A2(n1832), .ZN(n1723) );
  XNOR2_X1 U1833 ( .A(n1723), .B(KEYINPUT90), .ZN(n1725) );
  NAND2_X1 U1834 ( .A1(n1947), .A2(G326), .ZN(n1724) );
  NAND2_X1 U1835 ( .A1(n1725), .A2(n1724), .ZN(n1736) );
  NAND2_X1 U1836 ( .A1(G322), .A2(n1956), .ZN(n1727) );
  NAND2_X1 U1837 ( .A1(G311), .A2(n1953), .ZN(n1726) );
  NAND2_X1 U1838 ( .A1(n1727), .A2(n1726), .ZN(n1728) );
  NOR2_X1 U1839 ( .A1(n1941), .A2(n1728), .ZN(n1734) );
  NAND2_X1 U1840 ( .A1(n1952), .A2(G317), .ZN(n1730) );
  NAND2_X1 U1841 ( .A1(G329), .A2(n1943), .ZN(n1729) );
  NAND2_X1 U1842 ( .A1(n1730), .A2(n1729), .ZN(n1732) );
  AND2_X1 U1843 ( .A1(n1860), .A2(G294), .ZN(n1731) );
  NOR2_X1 U1844 ( .A1(n1732), .A2(n1731), .ZN(n1733) );
  NAND2_X1 U1845 ( .A1(n1734), .A2(n1733), .ZN(n1735) );
  NOR2_X1 U1846 ( .A1(n1736), .A2(n1735), .ZN(n1737) );
  NAND2_X1 U1847 ( .A1(n1738), .A2(n1737), .ZN(n1779) );
  NAND2_X1 U1848 ( .A1(n1022), .A2(n1739), .ZN(n1740) );
  XNOR2_X1 U1849 ( .A(n1740), .B(KEYINPUT62), .ZN(n1755) );
  NAND2_X1 U1850 ( .A1(G355), .A2(n1902), .ZN(n1752) );
  NOR2_X1 U1851 ( .A1(n1741), .A2(G116), .ZN(n1742) );
  XNOR2_X1 U1852 ( .A(n1742), .B(KEYINPUT60), .ZN(n1750) );
  XNOR2_X1 U1853 ( .A(G77), .B(G50), .ZN(n1744) );
  XNOR2_X1 U1854 ( .A(n1744), .B(n1743), .ZN(n2068) );
  NAND2_X1 U1855 ( .A1(G45), .A2(n2068), .ZN(n1747) );
  NOR2_X1 U1856 ( .A1(n2064), .A2(n2063), .ZN(n2030) );
  NAND2_X1 U1857 ( .A1(n2030), .A2(n1745), .ZN(n1746) );
  NAND2_X1 U1858 ( .A1(n1747), .A2(n1746), .ZN(n1748) );
  NOR2_X1 U1859 ( .A1(n1748), .A2(n1826), .ZN(n1749) );
  NOR2_X1 U1860 ( .A1(n1750), .A2(n1749), .ZN(n1751) );
  NAND2_X1 U1861 ( .A1(n1752), .A2(n1751), .ZN(n1753) );
  NAND2_X1 U1862 ( .A1(n1753), .A2(n1823), .ZN(n1754) );
  NAND2_X1 U1863 ( .A1(n1755), .A2(n1754), .ZN(n1775) );
  NAND2_X1 U1864 ( .A1(G58), .A2(n1956), .ZN(n1757) );
  NAND2_X1 U1865 ( .A1(n1757), .A2(n1756), .ZN(n1758) );
  XNOR2_X1 U1866 ( .A(n1758), .B(KEYINPUT86), .ZN(n1770) );
  NAND2_X1 U1867 ( .A1(G159), .A2(n1943), .ZN(n1760) );
  NAND2_X1 U1868 ( .A1(n1952), .A2(G68), .ZN(n1759) );
  NAND2_X1 U1869 ( .A1(n1760), .A2(n1759), .ZN(n1763) );
  NAND2_X1 U1870 ( .A1(G77), .A2(n1953), .ZN(n1761) );
  XNOR2_X1 U1871 ( .A(KEYINPUT87), .B(n1761), .ZN(n1762) );
  NOR2_X1 U1872 ( .A1(n1763), .A2(n1762), .ZN(n1764) );
  NAND2_X1 U1873 ( .A1(G97), .A2(n1860), .ZN(n1884) );
  NAND2_X1 U1874 ( .A1(n1764), .A2(n1884), .ZN(n1765) );
  XNOR2_X1 U1875 ( .A(KEYINPUT88), .B(n1765), .ZN(n1766) );
  XNOR2_X1 U1876 ( .A(n1766), .B(KEYINPUT61), .ZN(n1768) );
  NAND2_X1 U1877 ( .A1(G50), .A2(n1947), .ZN(n1767) );
  NAND2_X1 U1878 ( .A1(n1768), .A2(n1767), .ZN(n1769) );
  NOR2_X1 U1879 ( .A1(n1770), .A2(n1769), .ZN(n1771) );
  NAND2_X1 U1880 ( .A1(n1771), .A2(n1931), .ZN(n1772) );
  NOR2_X1 U1881 ( .A1(n1773), .A2(n1772), .ZN(n1774) );
  NOR2_X1 U1882 ( .A1(n1775), .A2(n1774), .ZN(n1776) );
  XNOR2_X1 U1883 ( .A(n1776), .B(KEYINPUT89), .ZN(n1777) );
  NOR2_X1 U1884 ( .A1(n1940), .A2(n1777), .ZN(n1778) );
  NAND2_X1 U1885 ( .A1(n1779), .A2(n1778), .ZN(n1780) );
  NAND2_X1 U1886 ( .A1(n1781), .A2(n1780), .ZN(G396) );
  NOR2_X1 U1887 ( .A1(n1783), .A2(n2021), .ZN(n1802) );
  BUF_X1 U1888 ( .A(n1784), .Z(n1785) );
  NAND2_X1 U1889 ( .A1(n1787), .A2(n1786), .ZN(n1788) );
  XNOR2_X1 U1890 ( .A(n1785), .B(n1788), .ZN(n1789) );
  NAND2_X1 U1891 ( .A1(n1789), .A2(n1796), .ZN(n1792) );
  OR2_X1 U1892 ( .A1(n1796), .A2(n1790), .ZN(n1791) );
  NAND2_X1 U1893 ( .A1(n1792), .A2(n1791), .ZN(n1794) );
  XOR2_X1 U1894 ( .A(KEYINPUT111), .B(KEYINPUT53), .Z(n1793) );
  XNOR2_X1 U1895 ( .A(n1794), .B(n1793), .ZN(n1800) );
  NOR2_X1 U1896 ( .A1(n1796), .A2(n1795), .ZN(n1797) );
  NAND2_X1 U1897 ( .A1(n1798), .A2(n1797), .ZN(n1799) );
  NAND2_X1 U1898 ( .A1(n1800), .A2(n1799), .ZN(n1801) );
  NAND2_X1 U1899 ( .A1(G283), .A2(n1953), .ZN(n1803) );
  NAND2_X1 U1900 ( .A1(n1804), .A2(n1803), .ZN(n1821) );
  NAND2_X1 U1901 ( .A1(G303), .A2(n1956), .ZN(n1806) );
  NAND2_X1 U1902 ( .A1(G116), .A2(n1946), .ZN(n1805) );
  NAND2_X1 U1903 ( .A1(n1806), .A2(n1805), .ZN(n1809) );
  NAND2_X1 U1904 ( .A1(G107), .A2(n1860), .ZN(n1807) );
  XNOR2_X1 U1905 ( .A(KEYINPUT113), .B(n1807), .ZN(n1808) );
  NOR2_X1 U1906 ( .A1(n1809), .A2(n1808), .ZN(n1818) );
  NAND2_X1 U1907 ( .A1(n1947), .A2(G311), .ZN(n1810) );
  XNOR2_X1 U1908 ( .A(n1810), .B(KEYINPUT54), .ZN(n1815) );
  NAND2_X1 U1909 ( .A1(G317), .A2(n1943), .ZN(n1812) );
  NAND2_X1 U1910 ( .A1(n1952), .A2(G294), .ZN(n1811) );
  NAND2_X1 U1911 ( .A1(n1812), .A2(n1811), .ZN(n1813) );
  NOR2_X1 U1912 ( .A1(n1941), .A2(n1813), .ZN(n1814) );
  NAND2_X1 U1913 ( .A1(n1815), .A2(n1814), .ZN(n1816) );
  XOR2_X1 U1914 ( .A(KEYINPUT114), .B(n1816), .Z(n1817) );
  NAND2_X1 U1915 ( .A1(n1818), .A2(n1817), .ZN(n1819) );
  XOR2_X1 U1916 ( .A(KEYINPUT115), .B(n1819), .Z(n1820) );
  NOR2_X1 U1917 ( .A1(n1821), .A2(n1820), .ZN(n1853) );
  NAND2_X1 U1918 ( .A1(G87), .A2(n1992), .ZN(n1822) );
  NAND2_X1 U1919 ( .A1(n1823), .A2(n1822), .ZN(n1828) );
  XOR2_X1 U1920 ( .A(G270), .B(G264), .Z(n1825) );
  XNOR2_X1 U1921 ( .A(G257), .B(G250), .ZN(n1824) );
  XNOR2_X1 U1922 ( .A(n1825), .B(n1824), .ZN(n2067) );
  NOR2_X1 U1923 ( .A1(n2067), .A2(n1826), .ZN(n1827) );
  NOR2_X1 U1924 ( .A1(n1828), .A2(n1827), .ZN(n1829) );
  NOR2_X1 U1925 ( .A1(n1940), .A2(n1829), .ZN(n1851) );
  NAND2_X1 U1926 ( .A1(n1946), .A2(G58), .ZN(n1830) );
  NAND2_X1 U1927 ( .A1(n1831), .A2(n1830), .ZN(n1845) );
  NAND2_X1 U1928 ( .A1(G77), .A2(n1832), .ZN(n1958) );
  NAND2_X1 U1929 ( .A1(n1956), .A2(G150), .ZN(n1833) );
  NAND2_X1 U1930 ( .A1(n1958), .A2(n1833), .ZN(n1842) );
  NAND2_X1 U1931 ( .A1(G137), .A2(n1943), .ZN(n1835) );
  NAND2_X1 U1932 ( .A1(G50), .A2(n1953), .ZN(n1834) );
  NAND2_X1 U1933 ( .A1(n1835), .A2(n1834), .ZN(n1838) );
  NAND2_X1 U1934 ( .A1(n1952), .A2(G159), .ZN(n1836) );
  NAND2_X1 U1935 ( .A1(n1931), .A2(n1836), .ZN(n1837) );
  NOR2_X1 U1936 ( .A1(n1838), .A2(n1837), .ZN(n1840) );
  NAND2_X1 U1937 ( .A1(n1947), .A2(G143), .ZN(n1839) );
  NAND2_X1 U1938 ( .A1(n1840), .A2(n1839), .ZN(n1841) );
  NOR2_X1 U1939 ( .A1(n1842), .A2(n1841), .ZN(n1843) );
  XOR2_X1 U1940 ( .A(KEYINPUT112), .B(n1843), .Z(n1844) );
  NOR2_X1 U1941 ( .A1(n1845), .A2(n1844), .ZN(n1849) );
  OR2_X1 U1942 ( .A1(n1846), .A2(n1785), .ZN(n1847) );
  XOR2_X1 U1943 ( .A(KEYINPUT116), .B(n1847), .Z(n1848) );
  NOR2_X1 U1944 ( .A1(n1849), .A2(n1848), .ZN(n1850) );
  NAND2_X1 U1945 ( .A1(n1851), .A2(n1850), .ZN(n1852) );
  NOR2_X1 U1946 ( .A1(n1853), .A2(n1852), .ZN(n1854) );
  XOR2_X1 U1947 ( .A(KEYINPUT117), .B(n1854), .Z(n1855) );
  XNOR2_X1 U1948 ( .A(n1903), .B(n2026), .ZN(n1858) );
  NOR2_X1 U1949 ( .A1(n1859), .A2(n1858), .ZN(n1912) );
  NAND2_X1 U1950 ( .A1(n1956), .A2(G143), .ZN(n1879) );
  NAND2_X1 U1951 ( .A1(G137), .A2(n1947), .ZN(n1867) );
  NAND2_X1 U1952 ( .A1(G50), .A2(n1946), .ZN(n1862) );
  NAND2_X1 U1953 ( .A1(G58), .A2(n1860), .ZN(n1861) );
  NAND2_X1 U1954 ( .A1(n1862), .A2(n1861), .ZN(n1865) );
  NAND2_X1 U1955 ( .A1(n1953), .A2(G159), .ZN(n1863) );
  XOR2_X1 U1956 ( .A(KEYINPUT122), .B(n1863), .Z(n1864) );
  NOR2_X1 U1957 ( .A1(n1865), .A2(n1864), .ZN(n1866) );
  NAND2_X1 U1958 ( .A1(n1867), .A2(n1866), .ZN(n1868) );
  XNOR2_X1 U1959 ( .A(n1868), .B(KEYINPUT20), .ZN(n1877) );
  NAND2_X1 U1960 ( .A1(n1943), .A2(G132), .ZN(n1869) );
  XNOR2_X1 U1961 ( .A(KEYINPUT19), .B(n1869), .ZN(n1872) );
  NAND2_X1 U1962 ( .A1(n1952), .A2(G150), .ZN(n1870) );
  NAND2_X1 U1963 ( .A1(n1931), .A2(n1870), .ZN(n1871) );
  NOR2_X1 U1964 ( .A1(n1872), .A2(n1871), .ZN(n1873) );
  XOR2_X1 U1965 ( .A(KEYINPUT121), .B(n1873), .Z(n1874) );
  NAND2_X1 U1966 ( .A1(n1875), .A2(n1874), .ZN(n1876) );
  NOR2_X1 U1967 ( .A1(n1877), .A2(n1876), .ZN(n1878) );
  NAND2_X1 U1968 ( .A1(n1879), .A2(n1878), .ZN(n1907) );
  NAND2_X1 U1969 ( .A1(n1943), .A2(G311), .ZN(n1881) );
  NAND2_X1 U1970 ( .A1(n1952), .A2(G283), .ZN(n1880) );
  NAND2_X1 U1971 ( .A1(n1881), .A2(n1880), .ZN(n1882) );
  NOR2_X1 U1972 ( .A1(n1883), .A2(n1882), .ZN(n1890) );
  NAND2_X1 U1973 ( .A1(n1885), .A2(n1884), .ZN(n1888) );
  NAND2_X1 U1974 ( .A1(G116), .A2(n1953), .ZN(n1886) );
  XNOR2_X1 U1975 ( .A(KEYINPUT21), .B(n1886), .ZN(n1887) );
  NOR2_X1 U1976 ( .A1(n1888), .A2(n1887), .ZN(n1889) );
  NAND2_X1 U1977 ( .A1(n1890), .A2(n1889), .ZN(n1901) );
  NAND2_X1 U1978 ( .A1(n1947), .A2(G303), .ZN(n1892) );
  NAND2_X1 U1979 ( .A1(n1956), .A2(G294), .ZN(n1891) );
  NAND2_X1 U1980 ( .A1(n1892), .A2(n1891), .ZN(n1893) );
  XOR2_X1 U1981 ( .A(KEYINPUT118), .B(n1893), .Z(n1895) );
  NAND2_X1 U1982 ( .A1(G107), .A2(n1946), .ZN(n1894) );
  NAND2_X1 U1983 ( .A1(n1895), .A2(n1894), .ZN(n1896) );
  XOR2_X1 U1984 ( .A(KEYINPUT119), .B(n1896), .Z(n1897) );
  NOR2_X1 U1985 ( .A1(n1898), .A2(n1897), .ZN(n1899) );
  XOR2_X1 U1986 ( .A(KEYINPUT120), .B(n1899), .Z(n1900) );
  NOR2_X1 U1987 ( .A1(n1901), .A2(n1900), .ZN(n1905) );
  AND2_X1 U1988 ( .A1(n1903), .A2(n1902), .ZN(n1904) );
  NOR2_X1 U1989 ( .A1(n1905), .A2(n1904), .ZN(n1906) );
  NAND2_X1 U1990 ( .A1(n1907), .A2(n1906), .ZN(n1909) );
  NOR2_X1 U1991 ( .A1(G77), .A2(n1965), .ZN(n1908) );
  NOR2_X1 U1992 ( .A1(n1909), .A2(n1908), .ZN(n1910) );
  NOR2_X1 U1993 ( .A1(n1940), .A2(n1910), .ZN(n1911) );
  INV_X1 U1994 ( .A(G213), .ZN(n1989) );
  NOR2_X1 U1995 ( .A1(G343), .A2(n1989), .ZN(n1914) );
  NAND2_X1 U1996 ( .A1(n1914), .A2(G2897), .ZN(n1915) );
  XNOR2_X1 U1997 ( .A(n1915), .B(KEYINPUT63), .ZN(n1916) );
  INV_X1 U1998 ( .A(KEYINPUT46), .ZN(n1917) );
  XNOR2_X1 U1999 ( .A(n1972), .B(n1917), .ZN(n1918) );
  XNOR2_X1 U2000 ( .A(n1919), .B(n1918), .ZN(n1920) );
  XNOR2_X1 U2001 ( .A(n1921), .B(KEYINPUT105), .ZN(n1977) );
  NAND2_X1 U2002 ( .A1(G159), .A2(n1946), .ZN(n1923) );
  NAND2_X1 U2003 ( .A1(G132), .A2(n1947), .ZN(n1922) );
  NAND2_X1 U2004 ( .A1(n1923), .A2(n1922), .ZN(n1938) );
  NAND2_X1 U2005 ( .A1(G137), .A2(n1956), .ZN(n1925) );
  NAND2_X1 U2006 ( .A1(G150), .A2(n1953), .ZN(n1924) );
  NAND2_X1 U2007 ( .A1(n1925), .A2(n1924), .ZN(n1929) );
  NAND2_X1 U2008 ( .A1(n1952), .A2(G143), .ZN(n1926) );
  NAND2_X1 U2009 ( .A1(n1927), .A2(n1926), .ZN(n1928) );
  NOR2_X1 U2010 ( .A1(n1929), .A2(n1928), .ZN(n1936) );
  NAND2_X1 U2011 ( .A1(n1943), .A2(G128), .ZN(n1930) );
  NAND2_X1 U2012 ( .A1(n1931), .A2(n1930), .ZN(n1934) );
  NOR2_X1 U2013 ( .A1(n1932), .A2(n2063), .ZN(n1933) );
  NOR2_X1 U2014 ( .A1(n1934), .A2(n1933), .ZN(n1935) );
  NAND2_X1 U2015 ( .A1(n1936), .A2(n1935), .ZN(n1937) );
  NOR2_X1 U2016 ( .A1(n1938), .A2(n1937), .ZN(n1939) );
  NOR2_X1 U2017 ( .A1(n1940), .A2(n1939), .ZN(n1964) );
  NOR2_X1 U2018 ( .A1(n1942), .A2(n1941), .ZN(n1945) );
  NAND2_X1 U2019 ( .A1(G303), .A2(n1943), .ZN(n1944) );
  NAND2_X1 U2020 ( .A1(n1945), .A2(n1944), .ZN(n1951) );
  NAND2_X1 U2021 ( .A1(n1946), .A2(G97), .ZN(n1949) );
  NAND2_X1 U2022 ( .A1(n1947), .A2(G294), .ZN(n1948) );
  NAND2_X1 U2023 ( .A1(n1949), .A2(n1948), .ZN(n1950) );
  NOR2_X1 U2024 ( .A1(n1951), .A2(n1950), .ZN(n1962) );
  NAND2_X1 U2025 ( .A1(n1952), .A2(G116), .ZN(n1955) );
  NAND2_X1 U2026 ( .A1(n1953), .A2(G107), .ZN(n1954) );
  NAND2_X1 U2027 ( .A1(n1955), .A2(n1954), .ZN(n1960) );
  NAND2_X1 U2028 ( .A1(G283), .A2(n1956), .ZN(n1957) );
  NAND2_X1 U2029 ( .A1(n1958), .A2(n1957), .ZN(n1959) );
  NOR2_X1 U2030 ( .A1(n1960), .A2(n1959), .ZN(n1961) );
  NAND2_X1 U2031 ( .A1(n1962), .A2(n1961), .ZN(n1963) );
  NAND2_X1 U2032 ( .A1(n1964), .A2(n1963), .ZN(n1967) );
  NOR2_X1 U2033 ( .A1(G68), .A2(n1965), .ZN(n1966) );
  NOR2_X1 U2034 ( .A1(n1967), .A2(n1966), .ZN(n1968) );
  XNOR2_X1 U2035 ( .A(n1968), .B(KEYINPUT45), .ZN(n1971) );
  NOR2_X1 U2036 ( .A1(n1969), .A2(n1516), .ZN(n1970) );
  NOR2_X1 U2037 ( .A1(n1971), .A2(n1970), .ZN(n1975) );
  AND2_X1 U2038 ( .A1(n1973), .A2(n1972), .ZN(n1974) );
  NOR2_X1 U2039 ( .A1(n1975), .A2(n1974), .ZN(n1976) );
  NAND2_X1 U2040 ( .A1(n1977), .A2(n1976), .ZN(G381) );
  NOR2_X1 U2041 ( .A1(G375), .A2(G378), .ZN(n1986) );
  NOR2_X1 U2042 ( .A1(G393), .A2(G396), .ZN(n1979) );
  XNOR2_X1 U2043 ( .A(n1979), .B(KEYINPUT124), .ZN(n1980) );
  NAND2_X1 U2044 ( .A1(n1981), .A2(n1980), .ZN(n1984) );
  XNOR2_X1 U2045 ( .A(KEYINPUT123), .B(n1982), .ZN(n1983) );
  NOR2_X1 U2046 ( .A1(n1984), .A2(n1983), .ZN(n1985) );
  INV_X1 U2047 ( .A(n1986), .ZN(n1987) );
  NOR2_X1 U2048 ( .A1(G343), .A2(n1987), .ZN(n1988) );
  NOR2_X1 U2049 ( .A1(n1989), .A2(n1988), .ZN(n1990) );
  NAND2_X1 U2050 ( .A1(G20), .A2(n1991), .ZN(n2050) );
  INV_X1 U2051 ( .A(n2050), .ZN(n2036) );
  NAND2_X1 U2052 ( .A1(n2036), .A2(n2030), .ZN(n1996) );
  NOR2_X1 U2053 ( .A1(G257), .A2(G264), .ZN(n1993) );
  NOR2_X1 U2054 ( .A1(n1993), .A2(n1992), .ZN(n1994) );
  NAND2_X1 U2055 ( .A1(n1994), .A2(G250), .ZN(n1995) );
  NAND2_X1 U2056 ( .A1(n1996), .A2(n1995), .ZN(n2015) );
  NAND2_X1 U2057 ( .A1(G270), .A2(G116), .ZN(n1998) );
  NAND2_X1 U2058 ( .A1(G97), .A2(G257), .ZN(n1997) );
  NAND2_X1 U2059 ( .A1(n1998), .A2(n1997), .ZN(n2001) );
  NAND2_X1 U2060 ( .A1(G264), .A2(G107), .ZN(n1999) );
  XOR2_X1 U2061 ( .A(KEYINPUT50), .B(n1999), .Z(n2000) );
  NOR2_X1 U2062 ( .A1(n2001), .A2(n2000), .ZN(n2003) );
  NAND2_X1 U2063 ( .A1(G250), .A2(G87), .ZN(n2002) );
  NAND2_X1 U2064 ( .A1(n2003), .A2(n2002), .ZN(n2012) );
  NAND2_X1 U2065 ( .A1(G232), .A2(G58), .ZN(n2005) );
  NAND2_X1 U2066 ( .A1(G68), .A2(G238), .ZN(n2004) );
  NAND2_X1 U2067 ( .A1(n2005), .A2(n2004), .ZN(n2009) );
  NAND2_X1 U2068 ( .A1(G226), .A2(G50), .ZN(n2007) );
  NAND2_X1 U2069 ( .A1(G77), .A2(G244), .ZN(n2006) );
  NAND2_X1 U2070 ( .A1(n2007), .A2(n2006), .ZN(n2008) );
  NOR2_X1 U2071 ( .A1(n2009), .A2(n2008), .ZN(n2010) );
  XNOR2_X1 U2072 ( .A(KEYINPUT49), .B(n2010), .ZN(n2011) );
  NOR2_X1 U2073 ( .A1(n2012), .A2(n2011), .ZN(n2013) );
  NOR2_X1 U2074 ( .A1(n1101), .A2(n2013), .ZN(n2014) );
  NOR2_X1 U2075 ( .A1(n2015), .A2(n2014), .ZN(G361) );
  INV_X1 U2076 ( .A(n2016), .ZN(n2017) );
  AND2_X1 U2077 ( .A1(n2018), .A2(n2017), .ZN(G372) );
  INV_X1 U2078 ( .A(n2019), .ZN(n2020) );
  NAND2_X1 U2079 ( .A1(n2021), .A2(n2020), .ZN(G399) );
  NAND2_X1 U2080 ( .A1(n2024), .A2(n2023), .ZN(n2025) );
  NOR2_X1 U2081 ( .A1(n2027), .A2(n2025), .ZN(n2029) );
  AND2_X1 U2082 ( .A1(n2027), .A2(n2026), .ZN(n2028) );
  NOR2_X1 U2083 ( .A1(n2029), .A2(n2028), .ZN(n2033) );
  NAND2_X1 U2084 ( .A1(n2031), .A2(n2030), .ZN(n2032) );
  NAND2_X1 U2085 ( .A1(n2033), .A2(n2032), .ZN(G364) );
  INV_X1 U2086 ( .A(G116), .ZN(n2035) );
  NOR2_X1 U2087 ( .A1(n2035), .A2(n2034), .ZN(n2037) );
  NAND2_X1 U2088 ( .A1(n2037), .A2(n2036), .ZN(n2038) );
  XNOR2_X1 U2089 ( .A(KEYINPUT126), .B(n2038), .ZN(n2062) );
  NOR2_X1 U2090 ( .A1(G13), .A2(n2027), .ZN(n2058) );
  INV_X1 U2091 ( .A(n2058), .ZN(n2052) );
  XOR2_X1 U2092 ( .A(n2040), .B(n2039), .Z(n2041) );
  NAND2_X1 U2093 ( .A1(n2041), .A2(G330), .ZN(n2048) );
  NAND2_X1 U2094 ( .A1(n2043), .A2(n2042), .ZN(n2044) );
  NAND2_X1 U2095 ( .A1(n2044), .A2(G369), .ZN(n2046) );
  XNOR2_X1 U2096 ( .A(n2046), .B(n2045), .ZN(n2047) );
  XNOR2_X1 U2097 ( .A(n2048), .B(n2047), .ZN(n2049) );
  NAND2_X1 U2098 ( .A1(n2050), .A2(n2049), .ZN(n2051) );
  NAND2_X1 U2099 ( .A1(n2052), .A2(n2051), .ZN(n2060) );
  NAND2_X1 U2100 ( .A1(G58), .A2(G50), .ZN(n2053) );
  XNOR2_X1 U2101 ( .A(n2053), .B(G68), .ZN(n2056) );
  NAND2_X1 U2102 ( .A1(n2054), .A2(G50), .ZN(n2055) );
  NAND2_X1 U2103 ( .A1(n2056), .A2(n2055), .ZN(n2057) );
  NAND2_X1 U2104 ( .A1(n2058), .A2(n2057), .ZN(n2059) );
  NAND2_X1 U2105 ( .A1(n2060), .A2(n2059), .ZN(n2061) );
  NAND2_X1 U2106 ( .A1(n2062), .A2(n2061), .ZN(G367) );
  NAND2_X1 U2107 ( .A1(n2064), .A2(n2063), .ZN(n2065) );
  NOR2_X1 U2108 ( .A1(G77), .A2(n2065), .ZN(G353) );
  XOR2_X1 U2109 ( .A(n2067), .B(n2066), .Z(G358) );
  XOR2_X1 U2110 ( .A(n2069), .B(n2068), .Z(G351) );
endmodule

