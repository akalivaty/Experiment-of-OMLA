//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n205), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(new_n229), .A2(new_n223), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n252), .B2(new_n201), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G159), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(G20), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT72), .B1(new_n262), .B2(KEYINPUT7), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT7), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT73), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n268), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n263), .A2(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n257), .B1(new_n273), .B2(new_n223), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n219), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n262), .A2(KEYINPUT7), .B1(new_n266), .B2(new_n270), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n256), .B1(new_n280), .B2(G68), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n281), .B2(KEYINPUT16), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n209), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(new_n210), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n278), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n285), .A2(new_n288), .B1(new_n287), .B2(new_n284), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT74), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(G226), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n266), .B(new_n294), .C1(G223), .C2(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G87), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(new_n292), .A3(G274), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n298), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n230), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n297), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n283), .A2(new_n290), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT17), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n283), .A2(KEYINPUT17), .A3(new_n290), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n303), .A2(G179), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n303), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n280), .A2(G68), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(KEYINPUT16), .A3(new_n257), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n278), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n274), .B2(new_n275), .ZN(new_n320));
  INV_X1    g0120(.A(new_n290), .ZN(new_n321));
  OAI211_X1 g0121(.A(KEYINPUT18), .B(new_n316), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n323), .A3(new_n326), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n313), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n292), .A2(G274), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n298), .ZN(new_n332));
  INV_X1    g0132(.A(new_n301), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(G226), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G222), .A2(G1698), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n293), .A2(G223), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n266), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(G77), .C2(new_n266), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(KEYINPUT66), .B2(new_n342), .C1(new_n304), .C2(new_n340), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n288), .B(G50), .C1(G1), .C2(new_n210), .ZN(new_n344));
  INV_X1    g0144(.A(new_n287), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(G50), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n284), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n210), .A2(G33), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n347), .A2(new_n349), .B1(G150), .B2(new_n254), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n203), .A2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n279), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT9), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n342), .A2(KEYINPUT66), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT66), .B(new_n342), .C1(new_n343), .C2(new_n354), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n340), .A2(new_n360), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n361), .B1(G169), .B2(new_n340), .C1(new_n352), .C2(new_n346), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n209), .B2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n288), .A2(new_n364), .B1(new_n363), .B2(new_n287), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n347), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OR3_X1    g0168(.A1(new_n368), .A2(KEYINPUT65), .A3(new_n348), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT65), .B1(new_n368), .B2(new_n348), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n278), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n266), .A2(G232), .A3(new_n293), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n206), .C2(new_n266), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n338), .ZN(new_n377));
  INV_X1    g0177(.A(G244), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n300), .B1(new_n378), .B2(new_n301), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n315), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n376), .B2(new_n338), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n360), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(G190), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n372), .C1(new_n304), .C2(new_n383), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n330), .A2(new_n359), .A3(new_n362), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n254), .A2(G50), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT69), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n348), .A2(new_n363), .B1(new_n210), .B2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n279), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT11), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT11), .ZN(new_n396));
  OR3_X1    g0196(.A1(new_n345), .A2(KEYINPUT12), .A3(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT12), .B1(new_n345), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n223), .B1(new_n209), .B2(G20), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n397), .A2(new_n398), .B1(new_n288), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT70), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G226), .A2(G1698), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n230), .B2(G1698), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n266), .B1(G33), .B2(G97), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n300), .B1(new_n405), .B2(new_n292), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n292), .A2(KEYINPUT67), .A3(new_n298), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT67), .B1(new_n292), .B2(new_n298), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n408), .A2(new_n409), .A3(new_n224), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  INV_X1    g0212(.A(new_n409), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(G238), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n230), .A2(G1698), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G226), .B2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n259), .A2(new_n261), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n416), .A2(new_n417), .B1(new_n258), .B2(new_n205), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n338), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n414), .A2(new_n419), .A3(new_n420), .A4(new_n300), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n411), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n419), .A3(new_n300), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(KEYINPUT68), .A3(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(G169), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n422), .A2(KEYINPUT14), .A3(G169), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n411), .A2(G179), .A3(new_n421), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n402), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n430), .ZN(new_n432));
  AOI211_X1 g0232(.A(KEYINPUT70), .B(new_n432), .C1(new_n427), .C2(new_n428), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n401), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n422), .A2(G200), .A3(new_n424), .ZN(new_n435));
  INV_X1    g0235(.A(new_n401), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n306), .B1(new_n423), .B2(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n421), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(new_n293), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n338), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n338), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n451), .A2(new_n450), .ZN(new_n453));
  INV_X1    g0253(.A(new_n331), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n452), .A2(G257), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(G169), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n263), .A2(new_n267), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n271), .A2(new_n272), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n206), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n254), .A2(G77), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT76), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT6), .ZN(new_n464));
  AND4_X1   g0264(.A1(G97), .A2(new_n462), .A3(new_n464), .A4(new_n206), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n462), .A2(new_n464), .B1(new_n207), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n460), .B1(new_n468), .B2(new_n210), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n278), .B1(new_n459), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n345), .A2(G97), .ZN(new_n471));
  AOI211_X1 g0271(.A(new_n278), .B(new_n287), .C1(new_n209), .C2(G33), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G97), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n456), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n448), .A2(new_n360), .A3(new_n455), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n448), .A2(new_n477), .A3(new_n360), .A4(new_n455), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n448), .A2(new_n455), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT77), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(G200), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n451), .A2(G274), .A3(new_n292), .A4(new_n450), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n451), .A2(new_n450), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n292), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(new_n231), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n338), .B2(new_n447), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n306), .B1(new_n482), .B2(new_n304), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n483), .A2(new_n490), .A3(new_n470), .A4(new_n473), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n207), .A2(G87), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n494));
  OAI211_X1 g0294(.A(G33), .B(G97), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(new_n210), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n259), .A2(new_n261), .A3(new_n210), .A4(G68), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n348), .A2(new_n205), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n278), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n368), .A2(new_n287), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n288), .B(G87), .C1(G1), .C2(new_n258), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n226), .B1(new_n209), .B2(G45), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n292), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT79), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n292), .A3(KEYINPUT79), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(new_n454), .B2(new_n450), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n259), .A2(new_n261), .A3(G238), .A4(new_n293), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n338), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n510), .A2(G190), .A3(new_n515), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n504), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n315), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n510), .A2(new_n360), .A3(new_n515), .ZN(new_n521));
  INV_X1    g0321(.A(new_n368), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n288), .B(new_n522), .C1(G1), .C2(new_n258), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n501), .A2(new_n502), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n480), .A2(new_n491), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n452), .A2(G270), .B1(new_n453), .B2(new_n454), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n266), .A2(G264), .A3(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n417), .A2(G303), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n259), .A2(new_n261), .A3(G257), .A4(new_n293), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n338), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n528), .A2(new_n533), .A3(G179), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n288), .B(G116), .C1(G1), .C2(new_n258), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n287), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n445), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(G20), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n278), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT20), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n535), .B(new_n537), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n528), .A2(new_n533), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n544), .A3(KEYINPUT21), .A4(G169), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n544), .A3(G169), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n544), .B1(G200), .B2(new_n546), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n306), .B2(new_n546), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n548), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n210), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n210), .A2(KEYINPUT81), .A3(G87), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT22), .B1(new_n417), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n562), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n266), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n561), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT24), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n559), .A2(new_n560), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n417), .A2(KEYINPUT22), .A3(new_n562), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n266), .B2(new_n564), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(KEYINPUT82), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n278), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n555), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n567), .A2(new_n568), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT24), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(KEYINPUT83), .A3(new_n278), .A4(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n472), .A2(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT25), .B1(new_n287), .B2(new_n206), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n417), .A2(new_n231), .A3(new_n293), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n259), .A2(new_n261), .A3(G250), .A4(new_n293), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n338), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n452), .A2(G264), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n484), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n306), .B2(new_n597), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n584), .A2(new_n590), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n589), .B1(new_n579), .B2(new_n583), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n315), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G179), .B2(new_n597), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n554), .B(new_n601), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  NOR4_X1   g0405(.A1(new_n389), .A2(new_n440), .A3(new_n527), .A4(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n385), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n439), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n313), .B1(new_n434), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n327), .A2(new_n322), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n359), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n362), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n389), .A2(new_n440), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n551), .A2(new_n545), .A3(new_n547), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n602), .B2(new_n604), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT84), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n589), .B(new_n599), .C1(new_n579), .C2(new_n583), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n527), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT84), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n615), .C1(new_n602), .C2(new_n604), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n474), .A2(new_n479), .A3(new_n525), .A4(new_n519), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n526), .A2(KEYINPUT26), .A3(new_n479), .A4(new_n474), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT85), .B1(new_n627), .B2(new_n525), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  INV_X1    g0429(.A(new_n525), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n625), .C2(new_n626), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n622), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n614), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n613), .A2(new_n633), .ZN(G369));
  INV_X1    g0434(.A(new_n554), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n544), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n615), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G330), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n604), .B1(new_n584), .B2(new_n590), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n618), .ZN(new_n651));
  INV_X1    g0451(.A(new_n641), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n602), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n650), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n644), .A2(new_n652), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n641), .B(KEYINPUT86), .Z(new_n659));
  AOI22_X1  g0459(.A1(new_n651), .A2(new_n658), .B1(new_n650), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n213), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n217), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n632), .A2(new_n659), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n480), .A2(new_n491), .A3(new_n526), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n616), .A2(new_n672), .A3(new_n601), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n627), .A2(new_n525), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n652), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT29), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(G179), .B1(new_n528), .B2(new_n533), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n481), .A3(new_n516), .A4(new_n597), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n515), .A2(new_n510), .A3(new_n595), .A4(new_n596), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n534), .A3(new_n488), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(KEYINPUT30), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n528), .A2(new_n533), .A3(G179), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n595), .A2(new_n596), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n516), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n687), .B2(new_n488), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n680), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n659), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  INV_X1    g0492(.A(new_n680), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n682), .A2(KEYINPUT30), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n687), .A2(new_n684), .A3(new_n488), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n692), .B1(new_n696), .B2(new_n652), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n651), .A2(new_n672), .A3(new_n554), .A4(new_n659), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n648), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n678), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n668), .B1(new_n704), .B2(G1), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT87), .Z(G364));
  NOR2_X1   g0506(.A1(new_n646), .A2(G330), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n286), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n209), .B1(new_n709), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n663), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n649), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n213), .A2(new_n266), .ZN(new_n715));
  INV_X1    g0515(.A(G355), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(G116), .B2(new_n213), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n662), .A2(new_n266), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n449), .B2(new_n218), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n247), .A2(new_n449), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n315), .A2(KEYINPUT89), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n210), .B1(KEYINPUT89), .B2(new_n315), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n219), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n712), .B1(new_n722), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n210), .A2(new_n360), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n304), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G317), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n210), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n734), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G303), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n740), .B1(new_n741), .B2(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n733), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n733), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n417), .B1(new_n747), .B2(new_n749), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  OR3_X1    g0554(.A1(KEYINPUT90), .A2(G179), .A3(G200), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT90), .B1(G179), .B2(G200), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n210), .B(G190), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n746), .B(new_n754), .C1(G329), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n306), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n210), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(new_n304), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n758), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT93), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n760), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G97), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n223), .B2(new_n735), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT91), .Z(new_n774));
  NAND2_X1  g0574(.A1(new_n757), .A2(G159), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT32), .Z(new_n776));
  OAI22_X1  g0576(.A1(new_n752), .A2(new_n229), .B1(new_n763), .B2(new_n202), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n266), .B1(new_n743), .B2(new_n206), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n225), .A2(new_n745), .B1(new_n749), .B2(new_n363), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n774), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n768), .A2(new_n769), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n770), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n732), .B1(new_n783), .B2(new_n726), .ZN(new_n784));
  INV_X1    g0584(.A(new_n729), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n646), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n714), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n373), .A2(new_n641), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n372), .B1(new_n315), .B2(new_n381), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n387), .A2(new_n789), .B1(new_n790), .B2(new_n384), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n385), .A2(new_n641), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT97), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT97), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n790), .A2(new_n384), .A3(new_n652), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n789), .A2(new_n387), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n607), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n669), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n798), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n632), .A2(new_n659), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n712), .B1(new_n802), .B2(new_n702), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n702), .B2(new_n802), .ZN(new_n804));
  INV_X1    g0604(.A(new_n726), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n728), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n712), .B1(new_n807), .B2(G77), .ZN(new_n808));
  INV_X1    g0608(.A(new_n749), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G150), .A2(new_n736), .B1(new_n809), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n763), .B2(new_n811), .C1(new_n812), .C2(new_n752), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n771), .A2(G58), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n266), .B1(new_n743), .B2(new_n223), .C1(new_n202), .C2(new_n745), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G132), .B2(new_n757), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n772), .B1(new_n761), .B2(new_n752), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT95), .Z(new_n822));
  OAI221_X1 g0622(.A(new_n417), .B1(new_n536), .B2(new_n749), .C1(new_n763), .C2(new_n744), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n743), .A2(new_n225), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n206), .A2(new_n745), .B1(new_n735), .B2(new_n741), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n757), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n747), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n820), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n808), .B1(new_n829), .B2(new_n726), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n800), .B2(new_n728), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n804), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n709), .A2(new_n209), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n429), .A2(new_n430), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT70), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n429), .A2(new_n402), .A3(new_n430), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n439), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n436), .A2(new_n652), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT99), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n839), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n434), .A2(new_n439), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n838), .A2(KEYINPUT99), .A3(new_n839), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n801), .A2(KEYINPUT98), .A3(new_n795), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT98), .B1(new_n801), .B2(new_n795), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT100), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  INV_X1    g0652(.A(new_n639), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n320), .B2(new_n321), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n325), .A2(new_n854), .A3(new_n855), .A4(new_n309), .ZN(new_n856));
  INV_X1    g0656(.A(new_n275), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n281), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n289), .B1(new_n319), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n289), .C1(new_n319), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n853), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n316), .A3(new_n862), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n863), .A2(new_n864), .A3(new_n309), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n856), .B1(new_n865), .B2(new_n855), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n330), .B2(new_n863), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n866), .B(KEYINPUT38), .C1(new_n330), .C2(new_n863), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n851), .A2(new_n852), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n325), .A2(new_n854), .A3(new_n309), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(new_n855), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n311), .A2(new_n312), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n854), .B1(new_n875), .B2(new_n610), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n868), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  MUX2_X1   g0678(.A(new_n878), .B(new_n871), .S(KEYINPUT39), .Z(new_n879));
  AOI21_X1  g0679(.A(new_n436), .B1(new_n836), .B2(new_n837), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n652), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n882), .B1(new_n611), .B2(new_n639), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n872), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n671), .A2(new_n614), .A3(new_n677), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n613), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n870), .A2(new_n877), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n889), .A2(new_n697), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n798), .B1(new_n700), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT99), .B1(new_n838), .B2(new_n839), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n845), .A2(new_n844), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n888), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT40), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT40), .B1(new_n869), .B2(new_n870), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n846), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n700), .A2(new_n890), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n614), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n902), .A2(new_n903), .A3(new_n648), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n834), .B1(new_n887), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n887), .B2(new_n905), .ZN(new_n907));
  INV_X1    g0707(.A(new_n468), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(KEYINPUT35), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(KEYINPUT35), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(G116), .A3(new_n220), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n217), .A2(new_n363), .A3(new_n252), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n223), .A2(G50), .ZN(new_n914));
  OAI211_X1 g0714(.A(G1), .B(new_n286), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(new_n912), .A3(new_n915), .ZN(G367));
  AND2_X1   g0716(.A1(new_n470), .A2(new_n473), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n480), .B(new_n491), .C1(new_n917), .C2(new_n659), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n474), .A2(new_n690), .A3(new_n479), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n651), .A2(new_n658), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n491), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n480), .B1(new_n654), .B2(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n921), .A2(KEYINPUT42), .B1(new_n923), .B2(new_n659), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT102), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(KEYINPUT42), .C2(new_n921), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n504), .A2(new_n652), .ZN(new_n929));
  MUX2_X1   g0729(.A(new_n526), .B(new_n630), .S(new_n929), .Z(new_n930));
  OR3_X1    g0730(.A1(new_n928), .A2(KEYINPUT43), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n930), .B(KEYINPUT43), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n656), .B1(new_n918), .B2(new_n919), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n660), .A2(new_n920), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT44), .Z(new_n941));
  INV_X1    g0741(.A(new_n656), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n660), .A2(new_n920), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT45), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n942), .B1(new_n941), .B2(new_n944), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n651), .A2(new_n658), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n655), .B2(new_n658), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(new_n649), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n703), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n663), .B(new_n952), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n710), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n939), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n731), .B1(new_n662), .B2(new_n522), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n718), .A2(new_n243), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n663), .B(new_n711), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n417), .B1(new_n749), .B2(new_n741), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n735), .A2(new_n761), .B1(new_n743), .B2(new_n205), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G317), .C2(new_n757), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n771), .A2(G107), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n745), .A2(new_n536), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT46), .Z(new_n964));
  AOI22_X1  g0764(.A1(new_n751), .A2(G303), .B1(new_n762), .B2(G311), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT106), .ZN(new_n967));
  INV_X1    g0767(.A(new_n745), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G58), .A2(new_n968), .B1(new_n736), .B2(G159), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n202), .B2(new_n749), .C1(new_n827), .C2(new_n811), .ZN(new_n970));
  INV_X1    g0770(.A(new_n743), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n417), .B1(new_n971), .B2(G77), .ZN(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n763), .B2(new_n812), .C1(new_n973), .C2(new_n752), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n760), .A2(new_n223), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n970), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n958), .B1(new_n785), .B2(new_n930), .C1(new_n978), .C2(new_n805), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n955), .A2(new_n979), .ZN(G387));
  NAND2_X1  g0780(.A1(new_n950), .A2(new_n711), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT107), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n655), .A2(new_n785), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n715), .A2(new_n665), .B1(G107), .B2(new_n213), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n665), .B(new_n449), .C1(new_n223), .C2(new_n363), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT50), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n284), .B2(G50), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n347), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n989), .A2(new_n719), .A3(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G45), .B2(new_n240), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT108), .B1(new_n989), .B2(new_n719), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n712), .B1(new_n993), .B2(new_n731), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n266), .B1(new_n743), .B2(new_n205), .C1(new_n752), .C2(new_n202), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G159), .B2(new_n762), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G77), .A2(new_n968), .B1(new_n736), .B2(new_n347), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n223), .B2(new_n749), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G150), .B2(new_n757), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n771), .A2(new_n522), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n266), .B1(new_n971), .B2(G116), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G303), .A2(new_n809), .B1(new_n736), .B2(G311), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n763), .B2(new_n753), .C1(new_n737), .C2(new_n752), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  OAI22_X1  g0805(.A1(new_n760), .A2(new_n741), .B1(new_n761), .B2(new_n745), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(KEYINPUT109), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT109), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1002), .B1(new_n764), .B2(new_n827), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n994), .B1(new_n1012), .B2(new_n726), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n982), .B1(new_n983), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n704), .A2(new_n950), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n664), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n704), .B2(new_n950), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(G393));
  AOI21_X1  g0819(.A(new_n664), .B1(new_n947), .B2(new_n1016), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT110), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n945), .A2(new_n1021), .A3(new_n946), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT110), .B(new_n942), .C1(new_n941), .C2(new_n944), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n1024), .B2(new_n1016), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n719), .A2(new_n250), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n730), .B1(new_n205), .B2(new_n213), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n712), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n771), .A2(G77), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n202), .B2(new_n735), .C1(new_n284), .C2(new_n749), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n751), .A2(G159), .B1(new_n762), .B2(G150), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT51), .Z(new_n1033));
  AOI211_X1 g0833(.A(new_n417), .B(new_n824), .C1(G68), .C2(new_n968), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n812), .C2(new_n827), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n827), .A2(new_n753), .B1(new_n741), .B2(new_n745), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n771), .A2(G116), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n761), .A2(new_n749), .B1(new_n735), .B2(new_n744), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n266), .B(new_n1040), .C1(G107), .C2(new_n971), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n751), .A2(G311), .B1(new_n762), .B2(G317), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1031), .A2(new_n1035), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1028), .B1(new_n1046), .B2(new_n726), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n920), .B2(new_n785), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1025), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n710), .B1(new_n1024), .B2(KEYINPUT111), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT111), .B2(new_n1024), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G390));
  AOI211_X1 g0853(.A(new_n648), .B(new_n798), .C1(new_n700), .C2(new_n890), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n893), .B2(new_n892), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n879), .B1(new_n849), .B2(new_n881), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n795), .B1(new_n675), .B2(new_n798), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n893), .B2(new_n892), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n882), .B1(new_n870), .B2(new_n877), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1056), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n701), .B(new_n800), .C1(new_n893), .C2(new_n892), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n1062), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n801), .A2(new_n795), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT98), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n801), .A2(KEYINPUT98), .A3(new_n795), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n882), .B1(new_n1074), .B2(new_n846), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1067), .B(new_n1069), .C1(new_n1075), .C2(new_n879), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n711), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n712), .B1(new_n807), .B2(new_n347), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1080));
  OR3_X1    g0880(.A1(new_n1080), .A2(new_n745), .A3(new_n973), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n745), .B2(new_n973), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n762), .A2(G128), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G132), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n266), .B1(new_n743), .B2(new_n202), .C1(new_n752), .C2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G125), .C2(new_n757), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n811), .A2(new_n735), .B1(new_n749), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n771), .B2(G159), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n417), .B1(new_n225), .B2(new_n745), .C1(new_n752), .C2(new_n536), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G283), .B2(new_n762), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n757), .A2(G294), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n735), .A2(new_n206), .B1(new_n743), .B2(new_n223), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G97), .B2(new_n809), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1029), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1099), .B2(new_n726), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n879), .B2(new_n728), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1078), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT116), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n605), .A2(new_n527), .A3(new_n690), .ZN(new_n1104));
  OAI211_X1 g0904(.A(G330), .B(new_n800), .C1(new_n1104), .C2(new_n698), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1055), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n847), .B2(new_n848), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1058), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1067), .B(new_n1109), .C1(new_n846), .C2(new_n1054), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n614), .A2(G330), .A3(new_n899), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n885), .A2(new_n613), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1103), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1113), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(KEYINPUT116), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT117), .B1(new_n1077), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1103), .B(new_n1113), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT116), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n664), .B1(new_n1077), .B2(new_n1118), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1102), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  AOI211_X1 g0929(.A(G41), .B(new_n266), .C1(new_n968), .C2(G77), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n206), .B2(new_n752), .C1(new_n536), .C2(new_n763), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G97), .A2(new_n736), .B1(new_n971), .B2(G58), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n368), .B2(new_n749), .C1(new_n827), .C2(new_n741), .ZN(new_n1133));
  OR3_X1    g0933(.A1(new_n1131), .A2(new_n1133), .A3(new_n975), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT58), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(G33), .A2(G41), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(G50), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n266), .B2(G41), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n809), .A2(G137), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n1085), .B2(new_n735), .C1(new_n745), .C2(new_n1088), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n751), .A2(G128), .B1(new_n762), .B2(G125), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n973), .C2(new_n760), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT120), .Z(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g0948(.A(G159), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT121), .B(G124), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1137), .B1(new_n1149), .B2(new_n743), .C1(new_n827), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1147), .B2(KEYINPUT59), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1141), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n712), .B1(G50), .B2(new_n807), .C1(new_n1153), .C2(new_n805), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n359), .A2(new_n362), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n353), .A2(new_n639), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1154), .B1(new_n1165), .B2(new_n727), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1163), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n893), .A2(new_n892), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n891), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n896), .B1(new_n894), .B2(KEYINPUT40), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1171), .B2(new_n648), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1163), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n898), .A2(G330), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n884), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n872), .A2(new_n883), .A3(new_n1174), .A4(new_n1172), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1166), .B1(new_n1178), .B2(new_n711), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1113), .B1(new_n1077), .B2(new_n1118), .ZN(new_n1180));
  AND4_X1   g0980(.A1(new_n872), .A2(new_n883), .A3(new_n1174), .A4(new_n1172), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n872), .A2(new_n883), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n663), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1066), .B(new_n1076), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1116), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1178), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1179), .B1(new_n1184), .B2(new_n1187), .ZN(G375));
  NOR2_X1   g0988(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1122), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n953), .B(KEYINPUT123), .Z(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT124), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1168), .A2(new_n727), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n712), .B1(new_n807), .B2(G68), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n266), .B1(new_n743), .B2(new_n229), .C1(new_n752), .C2(new_n811), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G132), .B2(new_n762), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n749), .A2(new_n973), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1149), .A2(new_n745), .B1(new_n735), .B2(new_n1088), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G128), .C2(new_n757), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(new_n202), .C2(new_n760), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n417), .B1(new_n743), .B2(new_n363), .C1(new_n752), .C2(new_n741), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G294), .B2(new_n762), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n757), .A2(G303), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n205), .A2(new_n745), .B1(new_n735), .B2(new_n536), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G107), .B2(new_n809), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1000), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1196), .B1(new_n1209), .B2(new_n726), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1115), .A2(new_n711), .B1(new_n1195), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1194), .A2(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G387), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n1052), .A3(new_n1050), .A4(new_n1215), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G378), .A2(G381), .A3(new_n1216), .A4(G375), .ZN(G407));
  INV_X1    g1017(.A(G375), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n640), .A3(new_n1128), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n663), .B1(new_n1189), .B2(KEYINPUT60), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1191), .B2(KEYINPUT60), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1212), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G384), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n832), .A3(new_n1212), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n640), .A2(G213), .A3(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1227), .B(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1192), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1186), .A2(new_n1178), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1179), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1124), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1127), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1102), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(G375), .B2(new_n1128), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n640), .A2(G213), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1221), .B1(new_n1229), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(G390), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(G393), .B(new_n787), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G387), .A2(new_n1052), .A3(new_n1050), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1238), .A2(new_n1239), .A3(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT125), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1238), .A2(new_n1227), .A3(new_n1253), .A4(new_n1239), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1249), .B(new_n1255), .C1(new_n1252), .C2(new_n1250), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT126), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1251), .A2(new_n1257), .A3(new_n1258), .A4(new_n1254), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1240), .A2(KEYINPUT62), .A3(new_n1227), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1251), .A2(new_n1258), .A3(new_n1254), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT126), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1241), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1256), .B1(new_n1264), .B2(new_n1247), .ZN(G405));
  XNOR2_X1  g1065(.A(G375), .B(new_n1128), .ZN(new_n1266));
  XOR2_X1   g1066(.A(new_n1266), .B(new_n1227), .Z(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1247), .ZN(G402));
endmodule


