

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603;

  XNOR2_X1 U328 ( .A(n461), .B(KEYINPUT45), .ZN(n462) );
  XNOR2_X1 U329 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n321) );
  XNOR2_X1 U331 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U332 ( .A(G50GAT), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U333 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U334 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U335 ( .A(n332), .B(n331), .ZN(n335) );
  XNOR2_X1 U336 ( .A(n423), .B(n388), .ZN(n392) );
  XNOR2_X1 U337 ( .A(n399), .B(n398), .ZN(n400) );
  NOR2_X1 U338 ( .A1(n489), .A2(n517), .ZN(n456) );
  XNOR2_X1 U339 ( .A(n337), .B(n424), .ZN(n481) );
  NOR2_X1 U340 ( .A1(n542), .A2(n483), .ZN(n579) );
  XNOR2_X1 U341 ( .A(n401), .B(n400), .ZN(n557) );
  INV_X1 U342 ( .A(G106GAT), .ZN(n457) );
  XNOR2_X1 U343 ( .A(KEYINPUT28), .B(n481), .ZN(n523) );
  XNOR2_X1 U344 ( .A(n485), .B(G183GAT), .ZN(n486) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U346 ( .A(n487), .B(n486), .ZN(G1350GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT89), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n315) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G155GAT), .Z(n299) );
  XNOR2_X1 U351 ( .A(G127GAT), .B(G148GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n301) );
  XNOR2_X1 U354 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U356 ( .A(n303), .B(n302), .Z(n313) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT2), .ZN(n328) );
  XOR2_X1 U359 ( .A(n328), .B(KEYINPUT4), .Z(n306) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n311) );
  XNOR2_X1 U362 ( .A(G134GAT), .B(G120GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n307), .B(KEYINPUT0), .ZN(n345) );
  XOR2_X1 U364 ( .A(G162GAT), .B(n345), .Z(n309) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G1GAT), .Z(n440) );
  XNOR2_X1 U366 ( .A(G29GAT), .B(n440), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(n315), .B(n314), .Z(n528) );
  XOR2_X1 U371 ( .A(KEYINPUT85), .B(KEYINPUT88), .Z(n317) );
  XNOR2_X1 U372 ( .A(G211GAT), .B(G204GAT), .ZN(n316) );
  XOR2_X1 U373 ( .A(n317), .B(n316), .Z(n319) );
  XOR2_X1 U374 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n318) );
  XOR2_X1 U375 ( .A(G22GAT), .B(G155GAT), .Z(n404) );
  XNOR2_X1 U376 ( .A(n387), .B(n404), .ZN(n320) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n323) );
  NAND2_X1 U378 ( .A1(n322), .A2(n323), .ZN(n327) );
  INV_X1 U379 ( .A(n322), .ZN(n325) );
  INV_X1 U380 ( .A(n323), .ZN(n324) );
  NAND2_X1 U381 ( .A1(n325), .A2(n324), .ZN(n326) );
  NAND2_X1 U382 ( .A1(n327), .A2(n326), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n328), .B(KEYINPUT22), .ZN(n330) );
  INV_X1 U384 ( .A(KEYINPUT23), .ZN(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n334) );
  XNOR2_X1 U386 ( .A(G197GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n353) );
  XNOR2_X1 U388 ( .A(n335), .B(n353), .ZN(n337) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(G78GAT), .ZN(n336) );
  XOR2_X1 U390 ( .A(n336), .B(G148GAT), .Z(n424) );
  XOR2_X1 U391 ( .A(G176GAT), .B(KEYINPUT20), .Z(n339) );
  XNOR2_X1 U392 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n352) );
  XOR2_X1 U394 ( .A(G71GAT), .B(G183GAT), .Z(n341) );
  NAND2_X1 U395 ( .A1(G227GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n344) );
  XOR2_X1 U397 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n343) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n354) );
  XOR2_X1 U400 ( .A(n344), .B(n354), .Z(n347) );
  XNOR2_X1 U401 ( .A(G113GAT), .B(n345), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n405) );
  XOR2_X1 U404 ( .A(n348), .B(n405), .Z(n350) );
  XNOR2_X1 U405 ( .A(G43GAT), .B(G190GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n536) );
  INV_X1 U408 ( .A(n536), .ZN(n542) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n368) );
  XOR2_X1 U410 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n360) );
  XOR2_X1 U411 ( .A(G92GAT), .B(KEYINPUT93), .Z(n356) );
  NAND2_X1 U412 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n357), .B(KEYINPUT76), .ZN(n395) );
  XNOR2_X1 U416 ( .A(n358), .B(n395), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n366) );
  XOR2_X1 U418 ( .A(KEYINPUT78), .B(G211GAT), .Z(n362) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(G183GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n418) );
  XOR2_X1 U421 ( .A(G64GAT), .B(KEYINPUT73), .Z(n364) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G204GAT), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n432) );
  XOR2_X1 U424 ( .A(n418), .B(n432), .Z(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U426 ( .A(n368), .B(n367), .Z(n530) );
  INV_X1 U427 ( .A(n530), .ZN(n510) );
  NOR2_X1 U428 ( .A1(n542), .A2(n510), .ZN(n369) );
  NOR2_X1 U429 ( .A1(n481), .A2(n369), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT25), .B(n370), .Z(n375) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n371) );
  XOR2_X1 U432 ( .A(n371), .B(n530), .Z(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n373) );
  NAND2_X1 U434 ( .A1(n481), .A2(n542), .ZN(n372) );
  XOR2_X1 U435 ( .A(n373), .B(n372), .Z(n562) );
  INV_X1 U436 ( .A(n562), .ZN(n584) );
  NOR2_X1 U437 ( .A1(n377), .A2(n584), .ZN(n374) );
  NOR2_X1 U438 ( .A1(n375), .A2(n374), .ZN(n376) );
  NOR2_X1 U439 ( .A1(n528), .A2(n376), .ZN(n382) );
  INV_X1 U440 ( .A(n523), .ZN(n378) );
  INV_X1 U441 ( .A(n528), .ZN(n507) );
  NOR2_X1 U442 ( .A1(n507), .A2(n377), .ZN(n534) );
  NAND2_X1 U443 ( .A1(n378), .A2(n534), .ZN(n539) );
  XNOR2_X1 U444 ( .A(n539), .B(KEYINPUT97), .ZN(n379) );
  AND2_X1 U445 ( .A1(n379), .A2(n542), .ZN(n380) );
  XNOR2_X1 U446 ( .A(KEYINPUT98), .B(n380), .ZN(n381) );
  NOR2_X1 U447 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U448 ( .A(n383), .B(KEYINPUT100), .Z(n496) );
  XOR2_X1 U449 ( .A(KEYINPUT72), .B(G92GAT), .Z(n385) );
  XNOR2_X1 U450 ( .A(G99GAT), .B(G85GAT), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n423) );
  AND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n386) );
  XOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n390) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(G106GAT), .ZN(n389) );
  XOR2_X1 U455 ( .A(n390), .B(n389), .Z(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n401) );
  XOR2_X1 U457 ( .A(G29GAT), .B(G43GAT), .Z(n394) );
  XNOR2_X1 U458 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n443) );
  XNOR2_X1 U460 ( .A(n443), .B(n395), .ZN(n399) );
  XOR2_X1 U461 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n397) );
  XNOR2_X1 U462 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(n557), .B(KEYINPUT36), .Z(n598) );
  NAND2_X1 U465 ( .A1(n496), .A2(n598), .ZN(n421) );
  XOR2_X1 U466 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n403) );
  XNOR2_X1 U467 ( .A(KEYINPUT82), .B(KEYINPUT80), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U469 ( .A(n404), .B(G78GAT), .Z(n407) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(n405), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U472 ( .A(n409), .B(n408), .Z(n411) );
  NAND2_X1 U473 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U475 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n413) );
  XNOR2_X1 U476 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U478 ( .A(n415), .B(n414), .Z(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n417) );
  XNOR2_X1 U480 ( .A(G71GAT), .B(G57GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n418), .B(n431), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n595) );
  NOR2_X1 U484 ( .A1(n421), .A2(n595), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n422), .B(KEYINPUT37), .ZN(n489) );
  XOR2_X1 U486 ( .A(n424), .B(n423), .Z(n436) );
  XOR2_X1 U487 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n426) );
  XNOR2_X1 U488 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U490 ( .A(KEYINPUT74), .B(G120GAT), .Z(n428) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U493 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U496 ( .A(n436), .B(n435), .Z(n488) );
  INV_X1 U497 ( .A(n488), .ZN(n591) );
  XOR2_X1 U498 ( .A(KEYINPUT41), .B(n591), .Z(n573) );
  XOR2_X1 U499 ( .A(G15GAT), .B(G197GAT), .Z(n438) );
  XNOR2_X1 U500 ( .A(G141GAT), .B(G22GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U502 ( .A(n439), .B(G36GAT), .Z(n442) );
  XNOR2_X1 U503 ( .A(n440), .B(G50GAT), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U505 ( .A(n443), .B(KEYINPUT65), .Z(n445) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U508 ( .A(n447), .B(n446), .Z(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n449) );
  XNOR2_X1 U510 ( .A(G169GAT), .B(G8GAT), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n451) );
  XNOR2_X1 U513 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U516 ( .A(n455), .B(n454), .Z(n546) );
  NAND2_X1 U517 ( .A1(n573), .A2(n546), .ZN(n517) );
  XOR2_X1 U518 ( .A(KEYINPUT105), .B(n456), .Z(n532) );
  NAND2_X1 U519 ( .A1(n532), .A2(n523), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n458) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(G1339GAT) );
  AND2_X1 U522 ( .A1(n595), .A2(n598), .ZN(n463) );
  INV_X1 U523 ( .A(KEYINPUT110), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n464), .A2(n591), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT111), .ZN(n466) );
  INV_X1 U526 ( .A(n546), .ZN(n587) );
  NOR2_X1 U527 ( .A1(n466), .A2(n587), .ZN(n476) );
  INV_X1 U528 ( .A(KEYINPUT47), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT107), .B(n595), .ZN(n554) );
  INV_X1 U530 ( .A(n557), .ZN(n578) );
  XOR2_X1 U531 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n468) );
  NAND2_X1 U532 ( .A1(n573), .A2(n587), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U534 ( .A1(n578), .A2(n469), .ZN(n470) );
  AND2_X1 U535 ( .A1(n554), .A2(n470), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n472), .B(n471), .ZN(n474) );
  INV_X1 U537 ( .A(KEYINPUT109), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U539 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n477), .B(KEYINPUT48), .ZN(n540) );
  NOR2_X1 U541 ( .A1(n540), .A2(n510), .ZN(n478) );
  XNOR2_X1 U542 ( .A(KEYINPUT54), .B(n478), .ZN(n479) );
  NAND2_X1 U543 ( .A1(n479), .A2(n507), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n480), .B(KEYINPUT64), .ZN(n585) );
  NOR2_X1 U545 ( .A1(n585), .A2(n481), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n482), .B(KEYINPUT55), .ZN(n483) );
  INV_X1 U547 ( .A(n579), .ZN(n484) );
  NOR2_X1 U548 ( .A1(n484), .A2(n554), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n485) );
  INV_X1 U550 ( .A(G50GAT), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n587), .A2(n488), .ZN(n498) );
  NOR2_X1 U552 ( .A1(n489), .A2(n498), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n490), .Z(n512) );
  NOR2_X1 U554 ( .A1(n512), .A2(n378), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT102), .B(n491), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1331GAT) );
  NAND2_X1 U557 ( .A1(n557), .A2(n595), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT16), .ZN(n495) );
  XNOR2_X1 U559 ( .A(KEYINPUT83), .B(n495), .ZN(n497) );
  NAND2_X1 U560 ( .A1(n497), .A2(n496), .ZN(n516) );
  NOR2_X1 U561 ( .A1(n498), .A2(n516), .ZN(n505) );
  NAND2_X1 U562 ( .A1(n505), .A2(n528), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT34), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n500), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n505), .A2(n530), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U568 ( .A1(n505), .A2(n536), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U570 ( .A(G15GAT), .B(n504), .Z(G1326GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n523), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U573 ( .A1(n512), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n512), .A2(n510), .ZN(n511) );
  XOR2_X1 U577 ( .A(G36GAT), .B(n511), .Z(G1329GAT) );
  INV_X1 U578 ( .A(KEYINPUT40), .ZN(n514) );
  NOR2_X1 U579 ( .A1(n512), .A2(n542), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n519) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n524), .A2(n528), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n530), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n536), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n526) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G78GAT), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n532), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  INV_X1 U601 ( .A(n534), .ZN(n535) );
  NOR2_X1 U602 ( .A1(n540), .A2(n535), .ZN(n561) );
  NAND2_X1 U603 ( .A1(n536), .A2(n561), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n378), .A2(n537), .ZN(n538) );
  NOR2_X1 U605 ( .A1(KEYINPUT112), .A2(n538), .ZN(n545) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U607 ( .A1(KEYINPUT112), .A2(n541), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n558) );
  NOR2_X1 U610 ( .A1(n558), .A2(n546), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(G1340GAT) );
  INV_X1 U613 ( .A(n573), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n549), .A2(n558), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n551) );
  XNOR2_X1 U616 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1341GAT) );
  NOR2_X1 U619 ( .A1(n558), .A2(n554), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT50), .B(n555), .Z(n556) );
  XNOR2_X1 U621 ( .A(G127GAT), .B(n556), .ZN(G1342GAT) );
  NOR2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(G1343GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT116), .B(n563), .Z(n570) );
  NAND2_X1 U627 ( .A1(n570), .A2(n587), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n566) );
  NAND2_X1 U630 ( .A1(n573), .A2(n570), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G148GAT), .B(n567), .ZN(G1345GAT) );
  XOR2_X1 U633 ( .A(G155GAT), .B(KEYINPUT117), .Z(n569) );
  NAND2_X1 U634 ( .A1(n595), .A2(n570), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n578), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n579), .A2(n587), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n575) );
  NAND2_X1 U642 ( .A1(n579), .A2(n573), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n581) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1351GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n589) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT123), .B(n586), .Z(n599) );
  NAND2_X1 U653 ( .A1(n599), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G197GAT), .B(n590), .ZN(G1352GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n593) );
  NAND2_X1 U657 ( .A1(n599), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(G204GAT), .B(n594), .ZN(G1353GAT) );
  XOR2_X1 U660 ( .A(G211GAT), .B(KEYINPUT125), .Z(n597) );
  NAND2_X1 U661 ( .A1(n599), .A2(n595), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n597), .B(n596), .ZN(G1354GAT) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n603) );
  XOR2_X1 U664 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n601) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U666 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U667 ( .A(n603), .B(n602), .ZN(G1355GAT) );
endmodule

