

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(n696), .A2(n595), .ZN(n663) );
  XNOR2_X1 U553 ( .A(KEYINPUT32), .B(KEYINPUT105), .ZN(n670) );
  XNOR2_X1 U554 ( .A(n671), .B(n670), .ZN(n725) );
  NOR2_X1 U555 ( .A1(G651), .A2(n572), .ZN(n799) );
  NOR2_X1 U556 ( .A1(n527), .A2(n526), .ZN(G164) );
  AND2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U558 ( .A1(G114), .A2(n889), .ZN(n520) );
  INV_X1 U559 ( .A(G2105), .ZN(n523) );
  AND2_X1 U560 ( .A1(n523), .A2(G2104), .ZN(n893) );
  NAND2_X1 U561 ( .A1(G102), .A2(n893), .ZN(n519) );
  NAND2_X1 U562 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n521), .Z(n894) );
  NAND2_X1 U565 ( .A1(G138), .A2(n894), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n522), .B(KEYINPUT94), .ZN(n525) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n523), .ZN(n890) );
  NAND2_X1 U568 ( .A1(n890), .A2(G126), .ZN(n524) );
  NAND2_X1 U569 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U570 ( .A1(G113), .A2(n889), .ZN(n529) );
  NAND2_X1 U571 ( .A1(G137), .A2(n894), .ZN(n528) );
  NAND2_X1 U572 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U573 ( .A(KEYINPUT66), .B(n530), .ZN(n536) );
  NAND2_X1 U574 ( .A1(G101), .A2(n893), .ZN(n531) );
  XNOR2_X1 U575 ( .A(n531), .B(KEYINPUT65), .ZN(n532) );
  XNOR2_X1 U576 ( .A(n532), .B(KEYINPUT23), .ZN(n534) );
  NAND2_X1 U577 ( .A1(G125), .A2(n890), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U579 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U580 ( .A(G651), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G543), .A2(n539), .ZN(n537) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n537), .Z(n797) );
  NAND2_X1 U583 ( .A1(n797), .A2(G64), .ZN(n538) );
  XNOR2_X1 U584 ( .A(n538), .B(KEYINPUT68), .ZN(n546) );
  XNOR2_X1 U585 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n544) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n572) );
  NOR2_X1 U587 ( .A1(n572), .A2(n539), .ZN(n793) );
  NAND2_X1 U588 ( .A1(G77), .A2(n793), .ZN(n542) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n540), .B(KEYINPUT64), .ZN(n794) );
  NAND2_X1 U591 ( .A1(G90), .A2(n794), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U593 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G52), .A2(n799), .ZN(n547) );
  XNOR2_X1 U596 ( .A(KEYINPUT69), .B(n547), .ZN(n548) );
  NOR2_X1 U597 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U598 ( .A1(n799), .A2(G51), .ZN(n550) );
  XOR2_X1 U599 ( .A(KEYINPUT79), .B(n550), .Z(n552) );
  NAND2_X1 U600 ( .A1(n797), .A2(G63), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n553), .ZN(n560) );
  NAND2_X1 U603 ( .A1(G89), .A2(n794), .ZN(n554) );
  XNOR2_X1 U604 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G76), .A2(n793), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U607 ( .A(KEYINPUT78), .B(n557), .Z(n558) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n558), .ZN(n559) );
  NOR2_X1 U609 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U610 ( .A(n561), .B(KEYINPUT7), .Z(n562) );
  XNOR2_X1 U611 ( .A(KEYINPUT80), .B(n562), .ZN(G168) );
  XOR2_X1 U612 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U613 ( .A1(n794), .A2(G88), .ZN(n563) );
  XNOR2_X1 U614 ( .A(n563), .B(KEYINPUT90), .ZN(n571) );
  NAND2_X1 U615 ( .A1(G62), .A2(n797), .ZN(n564) );
  XNOR2_X1 U616 ( .A(n564), .B(KEYINPUT88), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n793), .A2(G75), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U619 ( .A1(G50), .A2(n799), .ZN(n567) );
  XNOR2_X1 U620 ( .A(KEYINPUT89), .B(n567), .ZN(n568) );
  NOR2_X1 U621 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U622 ( .A1(n571), .A2(n570), .ZN(G303) );
  NAND2_X1 U623 ( .A1(n572), .A2(G87), .ZN(n577) );
  NAND2_X1 U624 ( .A1(G49), .A2(n799), .ZN(n574) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U626 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U627 ( .A1(n797), .A2(n575), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U629 ( .A(KEYINPUT85), .B(n578), .Z(G288) );
  NAND2_X1 U630 ( .A1(n793), .A2(G73), .ZN(n580) );
  XNOR2_X1 U631 ( .A(KEYINPUT2), .B(KEYINPUT86), .ZN(n579) );
  XNOR2_X1 U632 ( .A(n580), .B(n579), .ZN(n587) );
  NAND2_X1 U633 ( .A1(n797), .A2(G61), .ZN(n582) );
  NAND2_X1 U634 ( .A1(G86), .A2(n794), .ZN(n581) );
  NAND2_X1 U635 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U636 ( .A1(G48), .A2(n799), .ZN(n583) );
  XNOR2_X1 U637 ( .A(KEYINPUT87), .B(n583), .ZN(n584) );
  NOR2_X1 U638 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U639 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U640 ( .A1(G72), .A2(n793), .ZN(n589) );
  NAND2_X1 U641 ( .A1(G85), .A2(n794), .ZN(n588) );
  NAND2_X1 U642 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U643 ( .A(KEYINPUT67), .B(n590), .ZN(n594) );
  NAND2_X1 U644 ( .A1(G60), .A2(n797), .ZN(n592) );
  NAND2_X1 U645 ( .A1(G47), .A2(n799), .ZN(n591) );
  AND2_X1 U646 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U647 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X1 U648 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NAND2_X1 U649 ( .A1(G160), .A2(G40), .ZN(n695) );
  INV_X1 U650 ( .A(n695), .ZN(n595) );
  INV_X1 U651 ( .A(KEYINPUT100), .ZN(n596) );
  XNOR2_X1 U652 ( .A(n663), .B(n596), .ZN(n647) );
  NAND2_X1 U653 ( .A1(G2067), .A2(n647), .ZN(n598) );
  NAND2_X1 U654 ( .A1(G1348), .A2(n663), .ZN(n597) );
  NAND2_X1 U655 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U656 ( .A(n599), .B(KEYINPUT102), .ZN(n624) );
  NAND2_X1 U657 ( .A1(G79), .A2(n793), .ZN(n601) );
  NAND2_X1 U658 ( .A1(G66), .A2(n797), .ZN(n600) );
  NAND2_X1 U659 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U660 ( .A1(n799), .A2(G54), .ZN(n603) );
  NAND2_X1 U661 ( .A1(G92), .A2(n794), .ZN(n602) );
  NAND2_X1 U662 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U663 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n606) );
  XNOR2_X1 U665 ( .A(n607), .B(n606), .ZN(n978) );
  NAND2_X1 U666 ( .A1(G56), .A2(n797), .ZN(n608) );
  XOR2_X1 U667 ( .A(KEYINPUT14), .B(n608), .Z(n615) );
  NAND2_X1 U668 ( .A1(n793), .A2(G68), .ZN(n609) );
  XNOR2_X1 U669 ( .A(KEYINPUT75), .B(n609), .ZN(n612) );
  NAND2_X1 U670 ( .A1(G81), .A2(n794), .ZN(n610) );
  XOR2_X1 U671 ( .A(KEYINPUT12), .B(n610), .Z(n611) );
  NOR2_X1 U672 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U673 ( .A(n613), .B(KEYINPUT13), .ZN(n614) );
  NOR2_X1 U674 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U675 ( .A1(n799), .A2(G43), .ZN(n616) );
  NAND2_X1 U676 ( .A1(n617), .A2(n616), .ZN(n987) );
  INV_X1 U677 ( .A(G1996), .ZN(n618) );
  NOR2_X1 U678 ( .A1(n663), .A2(n618), .ZN(n619) );
  XOR2_X1 U679 ( .A(n619), .B(KEYINPUT26), .Z(n621) );
  NAND2_X1 U680 ( .A1(n663), .A2(G1341), .ZN(n620) );
  NAND2_X1 U681 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U682 ( .A1(n987), .A2(n622), .ZN(n634) );
  NOR2_X1 U683 ( .A1(n978), .A2(n634), .ZN(n623) );
  NOR2_X1 U684 ( .A1(n624), .A2(n623), .ZN(n638) );
  NAND2_X1 U685 ( .A1(G2072), .A2(n647), .ZN(n625) );
  XNOR2_X1 U686 ( .A(n625), .B(KEYINPUT27), .ZN(n627) );
  INV_X1 U687 ( .A(G1956), .ZN(n994) );
  NOR2_X1 U688 ( .A1(n647), .A2(n994), .ZN(n626) );
  NOR2_X1 U689 ( .A1(n627), .A2(n626), .ZN(n640) );
  NAND2_X1 U690 ( .A1(G65), .A2(n797), .ZN(n629) );
  NAND2_X1 U691 ( .A1(G53), .A2(n799), .ZN(n628) );
  NAND2_X1 U692 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U693 ( .A1(G78), .A2(n793), .ZN(n631) );
  NAND2_X1 U694 ( .A1(G91), .A2(n794), .ZN(n630) );
  NAND2_X1 U695 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U696 ( .A1(n633), .A2(n632), .ZN(n975) );
  NAND2_X1 U697 ( .A1(n640), .A2(n975), .ZN(n636) );
  NAND2_X1 U698 ( .A1(n634), .A2(n978), .ZN(n635) );
  NAND2_X1 U699 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U700 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U701 ( .A(KEYINPUT103), .B(n639), .Z(n643) );
  NOR2_X1 U702 ( .A1(n975), .A2(n640), .ZN(n641) );
  XNOR2_X1 U703 ( .A(KEYINPUT28), .B(n641), .ZN(n642) );
  NOR2_X1 U704 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U705 ( .A(n644), .B(KEYINPUT29), .ZN(n652) );
  INV_X1 U706 ( .A(n663), .ZN(n645) );
  NOR2_X1 U707 ( .A1(n645), .A2(G1961), .ZN(n646) );
  XNOR2_X1 U708 ( .A(n646), .B(KEYINPUT99), .ZN(n649) );
  XNOR2_X1 U709 ( .A(G2078), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U710 ( .A1(n647), .A2(n952), .ZN(n648) );
  NAND2_X1 U711 ( .A1(n649), .A2(n648), .ZN(n656) );
  NAND2_X1 U712 ( .A1(G171), .A2(n656), .ZN(n650) );
  XOR2_X1 U713 ( .A(KEYINPUT101), .B(n650), .Z(n651) );
  NAND2_X1 U714 ( .A1(n652), .A2(n651), .ZN(n661) );
  NAND2_X1 U715 ( .A1(G8), .A2(n663), .ZN(n731) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n731), .ZN(n677) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n663), .ZN(n672) );
  NOR2_X1 U718 ( .A1(n677), .A2(n672), .ZN(n653) );
  NAND2_X1 U719 ( .A1(G8), .A2(n653), .ZN(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U721 ( .A1(G168), .A2(n655), .ZN(n658) );
  NOR2_X1 U722 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U724 ( .A(KEYINPUT31), .B(n659), .Z(n660) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n674) );
  NAND2_X1 U726 ( .A1(n674), .A2(G286), .ZN(n662) );
  XNOR2_X1 U727 ( .A(n662), .B(KEYINPUT104), .ZN(n668) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n731), .ZN(n665) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n666), .A2(G303), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n669), .A2(G8), .ZN(n671) );
  NAND2_X1 U734 ( .A1(G8), .A2(n672), .ZN(n673) );
  XNOR2_X1 U735 ( .A(n673), .B(KEYINPUT98), .ZN(n675) );
  NAND2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U737 ( .A1(n677), .A2(n676), .ZN(n723) );
  INV_X1 U738 ( .A(n731), .ZN(n678) );
  NAND2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n969) );
  AND2_X1 U740 ( .A1(n678), .A2(n969), .ZN(n679) );
  NOR2_X1 U741 ( .A1(KEYINPUT33), .A2(n679), .ZN(n682) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NAND2_X1 U743 ( .A1(n977), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n680), .A2(n731), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n713) );
  XNOR2_X1 U746 ( .A(G1981), .B(KEYINPUT107), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n683), .B(G305), .ZN(n972) );
  XNOR2_X1 U748 ( .A(G2067), .B(KEYINPUT37), .ZN(n750) );
  NAND2_X1 U749 ( .A1(G104), .A2(n893), .ZN(n685) );
  NAND2_X1 U750 ( .A1(G140), .A2(n894), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n687) );
  XOR2_X1 U752 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n686) );
  XNOR2_X1 U753 ( .A(n687), .B(n686), .ZN(n692) );
  NAND2_X1 U754 ( .A1(G116), .A2(n889), .ZN(n689) );
  NAND2_X1 U755 ( .A1(G128), .A2(n890), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U757 ( .A(KEYINPUT35), .B(n690), .Z(n691) );
  NOR2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U759 ( .A(KEYINPUT36), .B(n693), .ZN(n880) );
  NOR2_X1 U760 ( .A1(n750), .A2(n880), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n694), .B(KEYINPUT96), .ZN(n938) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n752) );
  NAND2_X1 U763 ( .A1(n938), .A2(n752), .ZN(n697) );
  XOR2_X1 U764 ( .A(KEYINPUT97), .B(n697), .Z(n748) );
  NAND2_X1 U765 ( .A1(G129), .A2(n890), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G141), .A2(n894), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n893), .A2(G105), .ZN(n700) );
  XOR2_X1 U769 ( .A(KEYINPUT38), .B(n700), .Z(n701) );
  NOR2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n889), .A2(G117), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n886) );
  AND2_X1 U773 ( .A1(n886), .A2(G1996), .ZN(n922) );
  NAND2_X1 U774 ( .A1(G95), .A2(n893), .ZN(n706) );
  NAND2_X1 U775 ( .A1(G131), .A2(n894), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U777 ( .A1(G107), .A2(n889), .ZN(n708) );
  NAND2_X1 U778 ( .A1(G119), .A2(n890), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n885) );
  INV_X1 U781 ( .A(G1991), .ZN(n944) );
  NOR2_X1 U782 ( .A1(n885), .A2(n944), .ZN(n920) );
  OR2_X1 U783 ( .A1(n922), .A2(n920), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n752), .A2(n711), .ZN(n742) );
  AND2_X1 U785 ( .A1(n748), .A2(n742), .ZN(n733) );
  AND2_X1 U786 ( .A1(n972), .A2(n733), .ZN(n712) );
  AND2_X1 U787 ( .A1(n713), .A2(n712), .ZN(n720) );
  INV_X1 U788 ( .A(n720), .ZN(n714) );
  OR2_X1 U789 ( .A1(n723), .A2(n714), .ZN(n715) );
  NOR2_X1 U790 ( .A1(n725), .A2(n715), .ZN(n722) );
  NOR2_X1 U791 ( .A1(G1971), .A2(G303), .ZN(n984) );
  XOR2_X1 U792 ( .A(n984), .B(KEYINPUT106), .Z(n717) );
  INV_X1 U793 ( .A(KEYINPUT33), .ZN(n716) );
  NAND2_X1 U794 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U795 ( .A1(n718), .A2(n977), .ZN(n719) );
  AND2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U797 ( .A1(n722), .A2(n721), .ZN(n739) );
  NAND2_X1 U798 ( .A1(n731), .A2(n733), .ZN(n728) );
  OR2_X1 U799 ( .A1(n723), .A2(n728), .ZN(n724) );
  NOR2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n737) );
  NOR2_X1 U801 ( .A1(G2090), .A2(G303), .ZN(n726) );
  NAND2_X1 U802 ( .A1(G8), .A2(n726), .ZN(n727) );
  OR2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n735) );
  NOR2_X1 U804 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XOR2_X1 U805 ( .A(n729), .B(KEYINPUT24), .Z(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U812 ( .A1(n971), .A2(n752), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n755) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n886), .ZN(n917) );
  INV_X1 U815 ( .A(n742), .ZN(n745) );
  AND2_X1 U816 ( .A1(n944), .A2(n885), .ZN(n921) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n921), .A2(n743), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n917), .A2(n746), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT39), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n880), .A2(n750), .ZN(n927) );
  NAND2_X1 U824 ( .A1(n751), .A2(n927), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U827 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U828 ( .A(G2454), .B(G2443), .ZN(n766) );
  XOR2_X1 U829 ( .A(KEYINPUT108), .B(G2430), .Z(n758) );
  XNOR2_X1 U830 ( .A(G2446), .B(KEYINPUT109), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n758), .B(n757), .ZN(n762) );
  XOR2_X1 U832 ( .A(G2451), .B(G2427), .Z(n760) );
  XNOR2_X1 U833 ( .A(G1341), .B(G1348), .ZN(n759) );
  XNOR2_X1 U834 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U835 ( .A(n762), .B(n761), .Z(n764) );
  XNOR2_X1 U836 ( .A(G2435), .B(G2438), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n767) );
  AND2_X1 U839 ( .A1(n767), .A2(G14), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  XOR2_X1 U843 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n769) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n769), .B(n768), .ZN(G223) );
  XOR2_X1 U846 ( .A(G223), .B(KEYINPUT74), .Z(n834) );
  NAND2_X1 U847 ( .A1(n834), .A2(G567), .ZN(n770) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n770), .Z(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n778) );
  OR2_X1 U850 ( .A1(n987), .A2(n778), .ZN(n771) );
  XNOR2_X1 U851 ( .A(KEYINPUT76), .B(n771), .ZN(G153) );
  INV_X1 U852 ( .A(G171), .ZN(G301) );
  NAND2_X1 U853 ( .A1(G868), .A2(G301), .ZN(n773) );
  OR2_X1 U854 ( .A1(n978), .A2(G868), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n773), .A2(n772), .ZN(G284) );
  XNOR2_X1 U856 ( .A(n975), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U857 ( .A(KEYINPUT81), .B(G868), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G286), .A2(n774), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n775), .B(KEYINPUT82), .ZN(n777) );
  NOR2_X1 U860 ( .A1(G299), .A2(G868), .ZN(n776) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n778), .A2(G559), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n779), .A2(n978), .ZN(n780) );
  XNOR2_X1 U864 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n987), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G868), .A2(n978), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G123), .A2(n890), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n889), .A2(G111), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G99), .A2(n893), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G135), .A2(n894), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n919) );
  XNOR2_X1 U877 ( .A(n919), .B(G2096), .ZN(n792) );
  INV_X1 U878 ( .A(G2100), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(G156) );
  NAND2_X1 U880 ( .A1(G80), .A2(n793), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G93), .A2(n794), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n803) );
  NAND2_X1 U883 ( .A1(n797), .A2(G67), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n798), .B(KEYINPUT84), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n815) );
  NAND2_X1 U888 ( .A1(G559), .A2(n978), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n804), .B(KEYINPUT83), .ZN(n813) );
  XOR2_X1 U890 ( .A(n813), .B(n987), .Z(n805) );
  NOR2_X1 U891 ( .A1(G860), .A2(n805), .ZN(n806) );
  XOR2_X1 U892 ( .A(n815), .B(n806), .Z(G145) );
  INV_X1 U893 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U894 ( .A(G166), .B(n987), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(G299), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n808), .B(G305), .ZN(n809) );
  XNOR2_X1 U897 ( .A(n809), .B(G288), .ZN(n810) );
  XOR2_X1 U898 ( .A(n815), .B(n810), .Z(n812) );
  XNOR2_X1 U899 ( .A(G290), .B(KEYINPUT19), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n812), .B(n811), .ZN(n905) );
  XNOR2_X1 U901 ( .A(n813), .B(n905), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n814), .A2(G868), .ZN(n818) );
  INV_X1 U903 ( .A(G868), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n818), .A2(n817), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n819) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n820), .ZN(n822) );
  XOR2_X1 U909 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n821) );
  XNOR2_X1 U910 ( .A(n822), .B(n821), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n823), .A2(G2072), .ZN(n824) );
  XNOR2_X1 U912 ( .A(n824), .B(KEYINPUT92), .ZN(G158) );
  XOR2_X1 U913 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XOR2_X1 U914 ( .A(KEYINPUT93), .B(G44), .Z(n825) );
  XNOR2_X1 U915 ( .A(KEYINPUT3), .B(n825), .ZN(G218) );
  NAND2_X1 U916 ( .A1(G108), .A2(G120), .ZN(n826) );
  NOR2_X1 U917 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G69), .A2(n827), .ZN(n839) );
  NAND2_X1 U919 ( .A1(G567), .A2(n839), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U922 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U923 ( .A1(G96), .A2(n830), .ZN(n840) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n840), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n841) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U927 ( .A1(n841), .A2(n833), .ZN(n838) );
  NAND2_X1 U928 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(n834), .A2(G2106), .ZN(n835) );
  XNOR2_X1 U930 ( .A(n835), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U932 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(KEYINPUT111), .B(n841), .ZN(G319) );
  XOR2_X1 U943 ( .A(G2100), .B(G2096), .Z(n843) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2090), .Z(n845) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1981), .B(G1966), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n861) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G2474), .Z(n853) );
  XNOR2_X1 U956 ( .A(G1986), .B(KEYINPUT112), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U958 ( .A(G1976), .B(G1971), .Z(n855) );
  XNOR2_X1 U959 ( .A(G1961), .B(G1956), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U961 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U962 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U965 ( .A1(n890), .A2(G124), .ZN(n862) );
  XNOR2_X1 U966 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U967 ( .A1(G136), .A2(n894), .ZN(n863) );
  NAND2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n865), .B(KEYINPUT115), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G112), .A2(n889), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n893), .A2(G100), .ZN(n868) );
  XOR2_X1 U973 ( .A(KEYINPUT116), .B(n868), .Z(n869) );
  NOR2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT117), .B(n871), .Z(G162) );
  NAND2_X1 U976 ( .A1(G103), .A2(n893), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G139), .A2(n894), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G115), .A2(n889), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G127), .A2(n890), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n929) );
  XOR2_X1 U984 ( .A(G164), .B(n929), .Z(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U987 ( .A(n919), .B(KEYINPUT118), .ZN(n881) );
  XNOR2_X1 U988 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U989 ( .A(n884), .B(n883), .Z(n888) );
  XOR2_X1 U990 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U991 ( .A(n888), .B(n887), .ZN(n901) );
  NAND2_X1 U992 ( .A1(G118), .A2(n889), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U995 ( .A1(G106), .A2(n893), .ZN(n896) );
  NAND2_X1 U996 ( .A1(G142), .A2(n894), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(KEYINPUT45), .B(n897), .Z(n898) );
  NOR2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G160), .B(G162), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(G286), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(G171), .B(n978), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n908), .ZN(n909) );
  XOR2_X1 U1008 ( .A(KEYINPUT119), .B(n909), .Z(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n911), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(KEYINPUT120), .B(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n918), .Z(n936) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1026 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n964) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n964), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1038 ( .A(G1996), .B(G32), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(n944), .B(G25), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT122), .ZN(n949) );
  XOR2_X1 U1044 ( .A(G2067), .B(KEYINPUT123), .Z(n947) );
  XNOR2_X1 U1045 ( .A(G26), .B(n947), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G27), .B(n952), .Z(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT124), .B(n958), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(G34), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT125), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G2084), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n964), .B(n963), .ZN(n966) );
  INV_X1 U1058 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n967), .ZN(n1022) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n991) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT57), .ZN(n986) );
  XNOR2_X1 U1068 ( .A(n975), .B(n994), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1070 ( .A(n978), .B(G1348), .Z(n980) );
  XOR2_X1 U1071 ( .A(G171), .B(G1961), .Z(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1341), .B(n987), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n1020) );
  INV_X1 U1080 ( .A(G16), .ZN(n1018) );
  XNOR2_X1 U1081 ( .A(G20), .B(n994), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1087 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT126), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT60), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G5), .B(G1961), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(n1015), .B(KEYINPUT127), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

