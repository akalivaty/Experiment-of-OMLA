

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774;

  NAND2_X2 U377 ( .A1(n635), .A2(n613), .ZN(n417) );
  NOR2_X1 U378 ( .A1(G237), .A2(G953), .ZN(n464) );
  XNOR2_X1 U379 ( .A(n571), .B(KEYINPUT32), .ZN(n572) );
  XNOR2_X1 U380 ( .A(n374), .B(n405), .ZN(n667) );
  NOR2_X2 U381 ( .A1(n603), .A2(n638), .ZN(n371) );
  AND2_X2 U382 ( .A1(n379), .A2(n429), .ZN(n378) );
  AND2_X1 U383 ( .A1(n359), .A2(n427), .ZN(n377) );
  XNOR2_X2 U384 ( .A(n759), .B(n522), .ZN(n692) );
  XNOR2_X2 U385 ( .A(n430), .B(KEYINPUT22), .ZN(n578) );
  NOR2_X2 U386 ( .A1(n683), .A2(n687), .ZN(n685) );
  OR2_X1 U387 ( .A1(n692), .A2(n409), .ZN(n408) );
  INV_X2 U388 ( .A(G122), .ZN(n424) );
  AND2_X2 U389 ( .A1(n382), .A2(n380), .ZN(n717) );
  NAND2_X1 U390 ( .A1(n383), .A2(n367), .ZN(n382) );
  NAND2_X1 U391 ( .A1(n389), .A2(n386), .ZN(n575) );
  AND2_X1 U392 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U393 ( .A1(n620), .A2(n734), .ZN(n623) );
  XNOR2_X1 U394 ( .A(n371), .B(n370), .ZN(n620) );
  NAND2_X1 U395 ( .A1(n385), .A2(n637), .ZN(n388) );
  OR2_X1 U396 ( .A1(n676), .A2(n651), .ZN(n631) );
  OR2_X1 U397 ( .A1(n557), .A2(n556), .ZN(n562) );
  NOR2_X2 U398 ( .A1(n610), .A2(n608), .ZN(n586) );
  NAND2_X2 U399 ( .A1(n411), .A2(n408), .ZN(n588) );
  AND2_X1 U400 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U401 ( .A1(n410), .A2(n483), .ZN(n409) );
  XNOR2_X1 U402 ( .A(n423), .B(G101), .ZN(n520) );
  XNOR2_X1 U403 ( .A(KEYINPUT3), .B(G113), .ZN(n423) );
  XNOR2_X1 U404 ( .A(KEYINPUT4), .B(G146), .ZN(n488) );
  INV_X1 U405 ( .A(n645), .ZN(n357) );
  INV_X2 U406 ( .A(G116), .ZN(n425) );
  XNOR2_X2 U407 ( .A(n424), .B(G104), .ZN(n457) );
  XNOR2_X2 U408 ( .A(n425), .B(G107), .ZN(n470) );
  BUF_X1 U409 ( .A(n683), .Z(n750) );
  OR2_X1 U410 ( .A1(n719), .A2(G902), .ZN(n497) );
  INV_X1 U411 ( .A(G134), .ZN(n476) );
  NOR2_X1 U412 ( .A1(n750), .A2(n381), .ZN(n690) );
  NAND2_X1 U413 ( .A1(n667), .A2(n360), .ZN(n381) );
  NAND2_X1 U414 ( .A1(n403), .A2(n399), .ZN(n432) );
  AND2_X1 U415 ( .A1(n433), .A2(n404), .ZN(n403) );
  AND2_X1 U416 ( .A1(n577), .A2(n576), .ZN(n358) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n436) );
  XNOR2_X1 U418 ( .A(KEYINPUT5), .B(G119), .ZN(n516) );
  INV_X1 U419 ( .A(KEYINPUT48), .ZN(n405) );
  XOR2_X1 U420 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n473) );
  XNOR2_X1 U421 ( .A(n362), .B(G140), .ZN(n758) );
  XNOR2_X1 U422 ( .A(n469), .B(n468), .ZN(n557) );
  XNOR2_X1 U423 ( .A(n457), .B(n470), .ZN(n373) );
  XNOR2_X1 U424 ( .A(n420), .B(n414), .ZN(n419) );
  INV_X1 U425 ( .A(G110), .ZN(n420) );
  INV_X1 U426 ( .A(G119), .ZN(n414) );
  XNOR2_X1 U427 ( .A(n419), .B(G128), .ZN(n502) );
  XNOR2_X1 U428 ( .A(n758), .B(G146), .ZN(n498) );
  XNOR2_X1 U429 ( .A(n686), .B(n384), .ZN(n383) );
  XNOR2_X1 U430 ( .A(G137), .B(G131), .ZN(n487) );
  XOR2_X1 U431 ( .A(G107), .B(G110), .Z(n492) );
  XNOR2_X1 U432 ( .A(G140), .B(G101), .ZN(n493) );
  XNOR2_X1 U433 ( .A(n748), .B(n451), .ZN(n706) );
  INV_X1 U434 ( .A(n388), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n587), .B(KEYINPUT98), .ZN(n638) );
  NAND2_X1 U436 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U437 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U438 ( .A(n673), .B(KEYINPUT80), .ZN(n372) );
  INV_X1 U439 ( .A(G237), .ZN(n441) );
  INV_X1 U440 ( .A(G128), .ZN(n445) );
  XOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n447) );
  NAND2_X1 U442 ( .A1(n358), .A2(n436), .ZN(n426) );
  XNOR2_X1 U443 ( .A(n588), .B(KEYINPUT105), .ZN(n624) );
  NAND2_X1 U444 ( .A1(n667), .A2(n439), .ZN(n668) );
  INV_X1 U445 ( .A(KEYINPUT39), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n485), .B(n484), .ZN(n532) );
  XNOR2_X1 U447 ( .A(n557), .B(KEYINPUT102), .ZN(n533) );
  XNOR2_X1 U448 ( .A(n421), .B(n419), .ZN(n418) );
  XNOR2_X1 U449 ( .A(n373), .B(n520), .ZN(n422) );
  XNOR2_X1 U450 ( .A(n442), .B(KEYINPUT75), .ZN(n421) );
  XNOR2_X1 U451 ( .A(n438), .B(n437), .ZN(n712) );
  XNOR2_X1 U452 ( .A(n498), .B(G137), .ZN(n437) );
  XNOR2_X1 U453 ( .A(n462), .B(n465), .ZN(n369) );
  INV_X1 U454 ( .A(n690), .ZN(n380) );
  XNOR2_X1 U455 ( .A(n759), .B(n496), .ZN(n719) );
  XNOR2_X1 U456 ( .A(n646), .B(KEYINPUT36), .ZN(n647) );
  NAND2_X1 U457 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n415), .B(KEYINPUT109), .ZN(n682) );
  NOR2_X1 U459 ( .A1(n638), .A2(n416), .ZN(n415) );
  OR2_X1 U460 ( .A1(n639), .A2(n640), .ZN(n416) );
  AND2_X1 U461 ( .A1(n533), .A2(n532), .ZN(n734) );
  AND2_X1 U462 ( .A1(n679), .A2(n678), .ZN(n680) );
  AND2_X1 U463 ( .A1(n428), .A2(n594), .ZN(n359) );
  AND2_X1 U464 ( .A1(n619), .A2(n666), .ZN(n360) );
  XNOR2_X1 U465 ( .A(n432), .B(n366), .ZN(n554) );
  XOR2_X1 U466 ( .A(n488), .B(n487), .Z(n361) );
  INV_X1 U467 ( .A(n611), .ZN(n433) );
  XOR2_X1 U468 ( .A(G125), .B(KEYINPUT10), .Z(n362) );
  AND2_X1 U469 ( .A1(n396), .A2(n559), .ZN(n363) );
  AND2_X1 U470 ( .A1(n586), .A2(n649), .ZN(n364) );
  AND2_X1 U471 ( .A1(n393), .A2(n387), .ZN(n365) );
  XNOR2_X1 U472 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n366) );
  OR2_X1 U473 ( .A1(n689), .A2(n688), .ZN(n367) );
  XNOR2_X1 U474 ( .A(n463), .B(n369), .ZN(n700) );
  XNOR2_X1 U475 ( .A(n422), .B(n418), .ZN(n748) );
  INV_X1 U476 ( .A(n594), .ZN(n435) );
  AND2_X1 U477 ( .A1(n435), .A2(n436), .ZN(n368) );
  XNOR2_X2 U478 ( .A(n454), .B(n453), .ZN(n635) );
  NOR2_X1 U479 ( .A1(n665), .A2(n664), .ZN(n407) );
  XNOR2_X1 U480 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U481 ( .A1(n376), .A2(n378), .ZN(n683) );
  NAND2_X1 U482 ( .A1(n406), .A2(n407), .ZN(n374) );
  NAND2_X1 U483 ( .A1(n772), .A2(n770), .ZN(n573) );
  XNOR2_X2 U484 ( .A(n568), .B(KEYINPUT106), .ZN(n772) );
  NOR2_X1 U485 ( .A1(n372), .A2(n690), .ZN(n674) );
  NAND2_X1 U486 ( .A1(n375), .A2(n435), .ZN(n379) );
  NAND2_X1 U487 ( .A1(n427), .A2(n428), .ZN(n375) );
  NAND2_X1 U488 ( .A1(n377), .A2(n426), .ZN(n376) );
  XNOR2_X2 U489 ( .A(n489), .B(n361), .ZN(n759) );
  XNOR2_X2 U490 ( .A(n477), .B(n476), .ZN(n489) );
  XNOR2_X2 U491 ( .A(n446), .B(n445), .ZN(n477) );
  NAND2_X1 U492 ( .A1(n717), .A2(G217), .ZN(n713) );
  INV_X1 U493 ( .A(KEYINPUT83), .ZN(n384) );
  NAND2_X1 U494 ( .A1(n590), .A2(n555), .ZN(n385) );
  NAND2_X1 U495 ( .A1(n397), .A2(n363), .ZN(n392) );
  INV_X1 U496 ( .A(n554), .ZN(n397) );
  NAND2_X1 U497 ( .A1(n395), .A2(n365), .ZN(n386) );
  NOR2_X1 U498 ( .A1(n388), .A2(n559), .ZN(n387) );
  NAND2_X1 U499 ( .A1(n391), .A2(n559), .ZN(n390) );
  NAND2_X1 U500 ( .A1(n393), .A2(n394), .ZN(n391) );
  NAND2_X1 U501 ( .A1(n554), .A2(n555), .ZN(n393) );
  NOR2_X1 U502 ( .A1(n590), .A2(n555), .ZN(n396) );
  NAND2_X1 U503 ( .A1(n398), .A2(n434), .ZN(n399) );
  NAND2_X1 U504 ( .A1(n649), .A2(n586), .ZN(n398) );
  XNOR2_X2 U505 ( .A(n585), .B(KEYINPUT1), .ZN(n649) );
  NAND2_X1 U506 ( .A1(n400), .A2(n649), .ZN(n404) );
  NOR2_X1 U507 ( .A1(n610), .A2(n401), .ZN(n400) );
  NAND2_X1 U508 ( .A1(n402), .A2(KEYINPUT107), .ZN(n401) );
  INV_X1 U509 ( .A(n608), .ZN(n402) );
  XNOR2_X1 U510 ( .A(n633), .B(n632), .ZN(n406) );
  NAND2_X1 U511 ( .A1(n692), .A2(n524), .ZN(n413) );
  INV_X1 U512 ( .A(n524), .ZN(n410) );
  NAND2_X1 U513 ( .A1(n524), .A2(G902), .ZN(n412) );
  XNOR2_X2 U514 ( .A(n509), .B(n508), .ZN(n610) );
  NAND2_X1 U515 ( .A1(n682), .A2(n641), .ZN(n643) );
  XNOR2_X2 U516 ( .A(n623), .B(n622), .ZN(n716) );
  OR2_X2 U517 ( .A1(n639), .A2(n602), .ZN(n603) );
  NOR2_X2 U518 ( .A1(n709), .A2(n747), .ZN(n711) );
  NOR2_X2 U519 ( .A1(n696), .A2(n747), .ZN(n699) );
  XNOR2_X1 U520 ( .A(n503), .B(n500), .ZN(n438) );
  NAND2_X1 U521 ( .A1(n653), .A2(n551), .ZN(n553) );
  XNOR2_X2 U522 ( .A(n417), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X2 U523 ( .A(n560), .B(KEYINPUT88), .ZN(n427) );
  AND2_X2 U524 ( .A1(n574), .A2(n593), .ZN(n428) );
  NAND2_X1 U525 ( .A1(n358), .A2(n368), .ZN(n429) );
  NAND2_X1 U526 ( .A1(n578), .A2(n564), .ZN(n566) );
  NOR2_X2 U527 ( .A1(n561), .A2(n431), .ZN(n430) );
  NAND2_X1 U528 ( .A1(n563), .A2(n402), .ZN(n431) );
  INV_X1 U529 ( .A(KEYINPUT107), .ZN(n434) );
  NOR2_X2 U530 ( .A1(n703), .A2(n747), .ZN(n704) );
  NOR2_X2 U531 ( .A1(n714), .A2(n747), .ZN(n715) );
  AND2_X1 U532 ( .A1(n666), .A2(n774), .ZN(n439) );
  AND2_X1 U533 ( .A1(n772), .A2(n770), .ZN(n576) );
  XNOR2_X1 U534 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U535 ( .A(KEYINPUT82), .ZN(n669) );
  INV_X1 U536 ( .A(KEYINPUT68), .ZN(n565) );
  INV_X1 U537 ( .A(KEYINPUT89), .ZN(n646) );
  XNOR2_X1 U538 ( .A(n467), .B(n466), .ZN(n468) );
  AND2_X1 U539 ( .A1(n762), .A2(n695), .ZN(n747) );
  NAND2_X1 U540 ( .A1(G237), .A2(G234), .ZN(n440) );
  XNOR2_X1 U541 ( .A(n440), .B(KEYINPUT14), .ZN(n547) );
  NAND2_X1 U542 ( .A1(G952), .A2(n547), .ZN(n544) );
  INV_X1 U543 ( .A(G902), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n483), .A2(n441), .ZN(n452) );
  NAND2_X1 U545 ( .A1(n452), .A2(G214), .ZN(n613) );
  XNOR2_X1 U546 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n442) );
  XOR2_X1 U547 ( .A(KEYINPUT18), .B(G125), .Z(n444) );
  XNOR2_X2 U548 ( .A(KEYINPUT64), .B(G953), .ZN(n762) );
  INV_X1 U549 ( .A(n762), .ZN(n471) );
  NAND2_X1 U550 ( .A1(G224), .A2(n471), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n444), .B(n443), .ZN(n450) );
  XNOR2_X2 U552 ( .A(KEYINPUT67), .B(G143), .ZN(n446) );
  XNOR2_X1 U553 ( .A(n447), .B(n488), .ZN(n448) );
  XNOR2_X1 U554 ( .A(n477), .B(n448), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U556 ( .A(G902), .B(KEYINPUT15), .ZN(n687) );
  NAND2_X1 U557 ( .A1(n706), .A2(n687), .ZN(n454) );
  AND2_X1 U558 ( .A1(n452), .A2(G210), .ZN(n453) );
  INV_X1 U559 ( .A(KEYINPUT38), .ZN(n455) );
  XNOR2_X1 U560 ( .A(n635), .B(n455), .ZN(n601) );
  NAND2_X1 U561 ( .A1(n613), .A2(n601), .ZN(n456) );
  XNOR2_X1 U562 ( .A(n456), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U563 ( .A(n498), .B(G113), .ZN(n463) );
  XOR2_X1 U564 ( .A(n457), .B(G143), .Z(n461) );
  XOR2_X1 U565 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n459) );
  XNOR2_X1 U566 ( .A(G131), .B(KEYINPUT12), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U568 ( .A(KEYINPUT76), .B(n464), .ZN(n517) );
  AND2_X1 U569 ( .A1(n517), .A2(G214), .ZN(n465) );
  NOR2_X1 U570 ( .A1(n700), .A2(G902), .ZN(n469) );
  XNOR2_X1 U571 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n467) );
  INV_X1 U572 ( .A(G475), .ZN(n466) );
  XOR2_X1 U573 ( .A(n470), .B(KEYINPUT103), .Z(n475) );
  NAND2_X1 U574 ( .A1(G234), .A2(n471), .ZN(n472) );
  XNOR2_X1 U575 ( .A(n473), .B(n472), .ZN(n499) );
  NAND2_X1 U576 ( .A1(G217), .A2(n499), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n474), .B(n475), .ZN(n482) );
  XOR2_X1 U578 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n479) );
  XNOR2_X1 U579 ( .A(G122), .B(KEYINPUT9), .ZN(n478) );
  XNOR2_X1 U580 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U581 ( .A(n489), .B(n480), .ZN(n481) );
  XNOR2_X1 U582 ( .A(n482), .B(n481), .ZN(n743) );
  NAND2_X1 U583 ( .A1(n743), .A2(n483), .ZN(n485) );
  INV_X1 U584 ( .A(G478), .ZN(n484) );
  INV_X1 U585 ( .A(n532), .ZN(n556) );
  NOR2_X1 U586 ( .A1(n535), .A2(n562), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n486), .B(KEYINPUT41), .ZN(n676) );
  INV_X1 U588 ( .A(G227), .ZN(n490) );
  OR2_X1 U589 ( .A1(n762), .A2(n490), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n492), .B(n491), .ZN(n495) );
  XNOR2_X1 U591 ( .A(n493), .B(G104), .ZN(n494) );
  XNOR2_X1 U592 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X2 U593 ( .A(n497), .B(G469), .ZN(n585) );
  NAND2_X1 U594 ( .A1(G221), .A2(n499), .ZN(n500) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U597 ( .A1(G902), .A2(n712), .ZN(n509) );
  NAND2_X1 U598 ( .A1(n687), .A2(G234), .ZN(n505) );
  XNOR2_X1 U599 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n504) );
  XNOR2_X1 U600 ( .A(n505), .B(n504), .ZN(n510) );
  NAND2_X1 U601 ( .A1(G217), .A2(n510), .ZN(n507) );
  INV_X1 U602 ( .A(KEYINPUT25), .ZN(n506) );
  XOR2_X1 U603 ( .A(KEYINPUT21), .B(KEYINPUT97), .Z(n512) );
  NAND2_X1 U604 ( .A1(G221), .A2(n510), .ZN(n511) );
  XNOR2_X1 U605 ( .A(n512), .B(n511), .ZN(n608) );
  NOR2_X1 U606 ( .A1(n649), .A2(n586), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n513), .B(KEYINPUT50), .ZN(n514) );
  XNOR2_X1 U608 ( .A(n514), .B(KEYINPUT119), .ZN(n527) );
  AND2_X1 U609 ( .A1(n610), .A2(n608), .ZN(n515) );
  XOR2_X1 U610 ( .A(KEYINPUT49), .B(n515), .Z(n525) );
  XNOR2_X1 U611 ( .A(n516), .B(G116), .ZN(n519) );
  NAND2_X1 U612 ( .A1(n517), .A2(G210), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n519), .B(n518), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U615 ( .A(KEYINPUT73), .ZN(n523) );
  XNOR2_X1 U616 ( .A(n523), .B(G472), .ZN(n524) );
  NOR2_X1 U617 ( .A1(n525), .A2(n588), .ZN(n526) );
  NAND2_X1 U618 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n588), .A2(n364), .ZN(n582) );
  NAND2_X1 U620 ( .A1(n528), .A2(n582), .ZN(n529) );
  XNOR2_X1 U621 ( .A(KEYINPUT51), .B(n529), .ZN(n530) );
  NOR2_X1 U622 ( .A1(n676), .A2(n530), .ZN(n541) );
  XNOR2_X1 U623 ( .A(n588), .B(KEYINPUT6), .ZN(n611) );
  NOR2_X1 U624 ( .A1(n601), .A2(n613), .ZN(n531) );
  NOR2_X1 U625 ( .A1(n562), .A2(n531), .ZN(n537) );
  INV_X1 U626 ( .A(n734), .ZN(n534) );
  OR2_X1 U627 ( .A1(n533), .A2(n532), .ZN(n604) );
  AND2_X1 U628 ( .A1(n534), .A2(n604), .ZN(n657) );
  NOR2_X1 U629 ( .A1(n535), .A2(n657), .ZN(n536) );
  NOR2_X1 U630 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n538), .B(KEYINPUT120), .ZN(n539) );
  NOR2_X1 U632 ( .A1(n554), .A2(n539), .ZN(n540) );
  NOR2_X1 U633 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n542), .B(KEYINPUT52), .ZN(n543) );
  NOR2_X1 U635 ( .A1(n544), .A2(n543), .ZN(n675) );
  NOR2_X1 U636 ( .A1(G953), .A2(n544), .ZN(n546) );
  INV_X1 U637 ( .A(KEYINPUT94), .ZN(n545) );
  XNOR2_X1 U638 ( .A(n546), .B(n545), .ZN(n600) );
  NAND2_X1 U639 ( .A1(G902), .A2(n547), .ZN(n597) );
  INV_X1 U640 ( .A(G898), .ZN(n548) );
  NAND2_X1 U641 ( .A1(n548), .A2(G953), .ZN(n749) );
  OR2_X1 U642 ( .A1(n597), .A2(n749), .ZN(n549) );
  NAND2_X1 U643 ( .A1(n600), .A2(n549), .ZN(n550) );
  XOR2_X1 U644 ( .A(KEYINPUT95), .B(n550), .Z(n551) );
  XOR2_X1 U645 ( .A(KEYINPUT91), .B(KEYINPUT0), .Z(n552) );
  XNOR2_X1 U646 ( .A(n553), .B(n552), .ZN(n561) );
  BUF_X1 U647 ( .A(n561), .Z(n590) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n555) );
  AND2_X1 U649 ( .A1(n557), .A2(n556), .ZN(n637) );
  XOR2_X1 U650 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n558) );
  XNOR2_X1 U651 ( .A(KEYINPUT77), .B(n558), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n575), .A2(KEYINPUT44), .ZN(n560) );
  INV_X1 U653 ( .A(n562), .ZN(n563) );
  INV_X1 U654 ( .A(n624), .ZN(n595) );
  NOR2_X1 U655 ( .A1(n595), .A2(n649), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n566), .B(n565), .ZN(n567) );
  NAND2_X1 U657 ( .A1(n567), .A2(n610), .ZN(n568) );
  AND2_X1 U658 ( .A1(n610), .A2(n649), .ZN(n569) );
  AND2_X1 U659 ( .A1(n611), .A2(n569), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n578), .A2(n570), .ZN(n571) );
  XNOR2_X2 U661 ( .A(KEYINPUT78), .B(n572), .ZN(n770) );
  NAND2_X1 U662 ( .A1(n573), .A2(KEYINPUT44), .ZN(n574) );
  INV_X1 U663 ( .A(n575), .ZN(n577) );
  AND2_X1 U664 ( .A1(n578), .A2(n611), .ZN(n580) );
  INV_X1 U665 ( .A(n610), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U667 ( .A1(n649), .A2(n581), .ZN(n723) );
  NOR2_X1 U668 ( .A1(n590), .A2(n582), .ZN(n584) );
  XNOR2_X1 U669 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n737) );
  OR2_X1 U671 ( .A1(n638), .A2(n588), .ZN(n589) );
  NOR2_X1 U672 ( .A1(n590), .A2(n589), .ZN(n725) );
  NOR2_X1 U673 ( .A1(n737), .A2(n725), .ZN(n591) );
  NOR2_X1 U674 ( .A1(n657), .A2(n591), .ZN(n592) );
  NOR2_X1 U675 ( .A1(n723), .A2(n592), .ZN(n593) );
  XNOR2_X1 U676 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n594) );
  NAND2_X1 U677 ( .A1(n595), .A2(n613), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT30), .ZN(n639) );
  NOR2_X1 U679 ( .A1(G900), .A2(n597), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n598), .A2(n762), .ZN(n599) );
  AND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n607) );
  INV_X1 U682 ( .A(n607), .ZN(n634) );
  NAND2_X1 U683 ( .A1(n601), .A2(n634), .ZN(n602) );
  INV_X1 U684 ( .A(n604), .ZN(n736) );
  NAND2_X1 U685 ( .A1(n620), .A2(n736), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT114), .ZN(n774) );
  NAND2_X1 U687 ( .A1(n774), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X1 U688 ( .A(KEYINPUT79), .B(n606), .ZN(n619) );
  NOR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n734), .A2(n433), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n625), .A2(n612), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n644) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(n644), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n649), .A2(n615), .ZN(n617) );
  INV_X1 U696 ( .A(KEYINPUT43), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n617), .B(n616), .ZN(n618) );
  INV_X1 U698 ( .A(n635), .ZN(n645) );
  AND2_X1 U699 ( .A1(n618), .A2(n645), .ZN(n742) );
  INV_X1 U700 ( .A(n742), .ZN(n666) );
  INV_X1 U701 ( .A(KEYINPUT111), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT40), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U704 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n628), .A2(n585), .ZN(n651) );
  INV_X1 U707 ( .A(KEYINPUT113), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT42), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(n681) );
  NAND2_X1 U710 ( .A1(n716), .A2(n681), .ZN(n633) );
  XNOR2_X1 U711 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n657), .A2(KEYINPUT47), .ZN(n641) );
  AND2_X1 U713 ( .A1(n357), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n640) );
  INV_X1 U715 ( .A(KEYINPUT81), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n665) );
  NOR2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n740) );
  INV_X1 U719 ( .A(n651), .ZN(n652) );
  AND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n732) );
  NOR2_X1 U721 ( .A1(KEYINPUT47), .A2(KEYINPUT69), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n732), .A2(n654), .ZN(n656) );
  NAND2_X1 U723 ( .A1(KEYINPUT47), .A2(KEYINPUT69), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n659) );
  INV_X1 U725 ( .A(n657), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n662) );
  INV_X1 U727 ( .A(n732), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n660), .A2(KEYINPUT47), .ZN(n661) );
  AND2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n740), .A2(n663), .ZN(n664) );
  XNOR2_X2 U731 ( .A(n668), .B(KEYINPUT85), .ZN(n684) );
  NOR2_X1 U732 ( .A1(n684), .A2(KEYINPUT2), .ZN(n670) );
  XNOR2_X1 U733 ( .A(n670), .B(n669), .ZN(n672) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U735 ( .A1(n750), .A2(n688), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U738 ( .A1(n676), .A2(n554), .ZN(n677) );
  NOR2_X1 U739 ( .A1(G953), .A2(n677), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n680), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U741 ( .A(n681), .B(G137), .ZN(G39) );
  XNOR2_X1 U742 ( .A(n682), .B(G143), .ZN(G45) );
  NAND2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n687), .B(KEYINPUT84), .ZN(n689) );
  NAND2_X1 U745 ( .A1(n717), .A2(G472), .ZN(n694) );
  XOR2_X1 U746 ( .A(KEYINPUT93), .B(KEYINPUT62), .Z(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n694), .B(n693), .ZN(n696) );
  INV_X1 U749 ( .A(G952), .ZN(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n697), .B(KEYINPUT90), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(G57) );
  NAND2_X1 U753 ( .A1(n717), .A2(G475), .ZN(n702) );
  XOR2_X1 U754 ( .A(n700), .B(KEYINPUT59), .Z(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n704), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U757 ( .A1(n717), .A2(G210), .ZN(n708) );
  XNOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U761 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n710) );
  XNOR2_X1 U762 ( .A(n711), .B(n710), .ZN(G51) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U765 ( .A(n716), .B(G131), .ZN(G33) );
  NAND2_X1 U766 ( .A1(n717), .A2(G469), .ZN(n721) );
  XOR2_X1 U767 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n722), .A2(n747), .ZN(G54) );
  XOR2_X1 U771 ( .A(G101), .B(n723), .Z(G3) );
  NAND2_X1 U772 ( .A1(n725), .A2(n734), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(G104), .ZN(G6) );
  XNOR2_X1 U774 ( .A(G107), .B(KEYINPUT26), .ZN(n729) );
  XOR2_X1 U775 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n727) );
  NAND2_X1 U776 ( .A1(n725), .A2(n736), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(G9) );
  NAND2_X1 U779 ( .A1(n732), .A2(n736), .ZN(n731) );
  XOR2_X1 U780 ( .A(G128), .B(KEYINPUT29), .Z(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(G30) );
  NAND2_X1 U782 ( .A1(n732), .A2(n734), .ZN(n733) );
  XNOR2_X1 U783 ( .A(G146), .B(n733), .ZN(G48) );
  NAND2_X1 U784 ( .A1(n737), .A2(n734), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n735), .B(G113), .ZN(G15) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(G116), .ZN(G18) );
  XOR2_X1 U788 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(G125), .B(n741), .ZN(G27) );
  XOR2_X1 U791 ( .A(G140), .B(n742), .Z(G42) );
  NAND2_X1 U792 ( .A1(n717), .A2(G478), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n743), .B(KEYINPUT121), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n747), .A2(n746), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n757) );
  OR2_X1 U797 ( .A1(G953), .A2(n750), .ZN(n754) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(KEYINPUT123), .ZN(n756) );
  XNOR2_X1 U803 ( .A(n757), .B(n756), .ZN(G69) );
  XNOR2_X1 U804 ( .A(n758), .B(n759), .ZN(n764) );
  XNOR2_X1 U805 ( .A(n764), .B(KEYINPUT124), .ZN(n760) );
  XNOR2_X1 U806 ( .A(n684), .B(n760), .ZN(n761) );
  NOR2_X1 U807 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n763), .B(KEYINPUT125), .ZN(n769) );
  XNOR2_X1 U809 ( .A(n764), .B(G227), .ZN(n765) );
  NAND2_X1 U810 ( .A1(n765), .A2(G900), .ZN(n766) );
  XNOR2_X1 U811 ( .A(KEYINPUT126), .B(n766), .ZN(n767) );
  NAND2_X1 U812 ( .A1(n767), .A2(G953), .ZN(n768) );
  NAND2_X1 U813 ( .A1(n769), .A2(n768), .ZN(G72) );
  XNOR2_X1 U814 ( .A(G119), .B(n770), .ZN(G21) );
  XNOR2_X1 U815 ( .A(G122), .B(KEYINPUT127), .ZN(n771) );
  XNOR2_X1 U816 ( .A(n771), .B(n575), .ZN(G24) );
  XOR2_X1 U817 ( .A(n772), .B(G110), .Z(n773) );
  XNOR2_X1 U818 ( .A(KEYINPUT117), .B(n773), .ZN(G12) );
  XNOR2_X1 U819 ( .A(G134), .B(n774), .ZN(G36) );
endmodule

