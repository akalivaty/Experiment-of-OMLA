//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  AND2_X1   g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  NOR4_X1   g0019(.A1(new_n214), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n204), .ZN(new_n232));
  INV_X1    g0032(.A(G68), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n209), .B(new_n230), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n216), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G179), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G87), .ZN(new_n254));
  OR2_X1    g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(G226), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G223), .A2(G1698), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT73), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n265), .A2(new_n266), .A3(new_n269), .A4(G232), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT74), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT64), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n273), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(G274), .A3(new_n275), .A4(new_n265), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n272), .B1(new_n271), .B2(new_n276), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n253), .B(new_n263), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n263), .B1(new_n277), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT75), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(KEYINPUT75), .B(new_n263), .C1(new_n277), .C2(new_n278), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n231), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n257), .B2(G20), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n233), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n234), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n226), .A2(new_n233), .ZN(new_n299));
  OAI21_X1  g0099(.A(G20), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G159), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n300), .B(KEYINPUT72), .C1(new_n301), .C2(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n290), .B1(new_n308), .B2(KEYINPUT16), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n297), .B2(new_n304), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n288), .B(new_n231), .C1(G1), .C2(new_n204), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n313), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT18), .B1(new_n287), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(G169), .B1(new_n283), .B2(new_n284), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n309), .B2(new_n311), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT18), .ZN(new_n324));
  NOR4_X1   g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n280), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n271), .A2(new_n276), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT75), .B1(new_n331), .B2(new_n263), .ZN(new_n332));
  INV_X1    g0132(.A(new_n284), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n286), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(new_n320), .A3(new_n279), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n326), .A3(new_n324), .ZN(new_n336));
  AOI21_X1  g0136(.A(G200), .B1(new_n283), .B2(new_n284), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n331), .A2(new_n338), .A3(new_n263), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n323), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT17), .B(new_n323), .C1(new_n337), .C2(new_n340), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n336), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n327), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n258), .A2(G222), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G223), .A2(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n257), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n262), .C1(G77), .C2(new_n257), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n265), .A2(new_n266), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n276), .C1(new_n222), .C2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(G179), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n317), .A2(new_n221), .ZN(new_n354));
  OAI21_X1  g0154(.A(G20), .B1(new_n234), .B2(G50), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n204), .A2(G33), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n355), .B1(new_n356), .B2(new_n303), .C1(new_n357), .C2(new_n313), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n358), .B2(new_n289), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G50), .B2(new_n314), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n352), .A2(new_n286), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n353), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT66), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n352), .A2(new_n338), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(G200), .B2(new_n352), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n360), .A2(new_n364), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT67), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n371), .B(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT10), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n371), .B(KEYINPUT67), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n367), .A4(new_n369), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n363), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n346), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT13), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n265), .A2(G238), .A3(new_n266), .ZN(new_n381));
  OAI211_X1 g0181(.A(G232), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(G226), .B(new_n258), .C1(new_n293), .C2(new_n294), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n257), .A2(KEYINPUT68), .A3(G226), .A4(new_n258), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n381), .B1(new_n390), .B2(new_n262), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n380), .B1(new_n391), .B2(new_n276), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n265), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  INV_X1    g0194(.A(new_n276), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n394), .A2(KEYINPUT13), .A3(new_n395), .A4(new_n381), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(G190), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n303), .A2(new_n221), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n357), .A2(new_n223), .B1(new_n204), .B2(G68), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n289), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n401), .A2(KEYINPUT11), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(KEYINPUT11), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n315), .A2(new_n233), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n317), .A2(new_n233), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT69), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT70), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT70), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n404), .A2(new_n411), .A3(new_n406), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(G200), .B1(new_n392), .B2(new_n396), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n398), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT71), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT71), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n398), .A2(new_n413), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(G169), .B1(new_n392), .B2(new_n396), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT14), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n393), .A2(G179), .A3(new_n397), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(G169), .C1(new_n392), .C2(new_n396), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n413), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n317), .A2(new_n223), .ZN(new_n428));
  INV_X1    g0228(.A(new_n313), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n302), .B1(G20), .B2(G77), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n357), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n433), .B2(new_n289), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n314), .A2(G77), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G238), .A2(G1698), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n257), .B(new_n438), .C1(new_n227), .C2(G1698), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n262), .C1(G107), .C2(new_n257), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n276), .C1(new_n224), .C2(new_n351), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n286), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT65), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n437), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(G179), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n437), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n441), .A2(new_n338), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(G200), .B2(new_n441), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n419), .A2(new_n427), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n379), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n203), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n314), .A2(new_n455), .A3(new_n231), .A4(new_n288), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n315), .A2(new_n215), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT77), .B(G97), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n204), .B(new_n460), .C1(new_n461), .C2(G33), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n288), .A2(new_n231), .B1(G20), .B2(new_n215), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT20), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n458), .B(new_n459), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G264), .A2(G1698), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n257), .B(new_n467), .C1(new_n213), .C2(G1698), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT82), .B(G303), .Z(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n262), .C1(new_n257), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n203), .A2(G45), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(G274), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n262), .B1(new_n474), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G270), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(G169), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(new_n253), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n466), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n466), .A2(new_n478), .A3(KEYINPUT21), .A4(G169), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n204), .A2(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT23), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  AOI21_X1  g0289(.A(G20), .B1(new_n255), .B2(new_n256), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G87), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n204), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(new_n488), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT24), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n492), .B(KEYINPUT22), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT24), .A3(new_n486), .A4(new_n488), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n498), .A3(new_n289), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n457), .A2(G107), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n314), .A2(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n476), .A2(G264), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n211), .A2(new_n258), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n257), .B(new_n505), .C1(G257), .C2(new_n258), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n265), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n475), .ZN(new_n509));
  NOR4_X1   g0309(.A1(new_n504), .A2(new_n508), .A3(new_n509), .A4(G179), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n286), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n485), .B1(new_n503), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n457), .A2(new_n431), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n461), .B2(new_n357), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n257), .A2(new_n204), .A3(G68), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G87), .A2(G107), .ZN(new_n518));
  AND2_X1   g0318(.A1(KEYINPUT77), .A2(G97), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT77), .A2(G97), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n204), .B1(new_n389), .B2(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n289), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n431), .A2(new_n314), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT81), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  AOI211_X1 g0329(.A(new_n529), .B(new_n526), .C1(new_n524), .C2(new_n289), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n514), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n224), .A2(G1698), .ZN(new_n533));
  OAI221_X1 g0333(.A(new_n533), .B1(G238), .B2(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n532), .A3(new_n535), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n262), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n473), .A2(new_n262), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n211), .B2(new_n472), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n253), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n286), .A3(new_n541), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n531), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(G68), .A2(new_n490), .B1(new_n521), .B2(new_n522), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n290), .B1(new_n546), .B2(new_n516), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n529), .B1(new_n547), .B2(new_n526), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n534), .A2(new_n532), .A3(new_n535), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n551), .A2(new_n536), .A3(new_n265), .ZN(new_n552));
  INV_X1    g0352(.A(new_n541), .ZN(new_n553));
  OAI21_X1  g0353(.A(G190), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n456), .A2(new_n210), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n539), .A2(G200), .A3(new_n541), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n550), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n545), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n511), .A2(new_n338), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n561));
  INV_X1    g0361(.A(G200), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n503), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n478), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n466), .B1(new_n566), .B2(G190), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(G244), .C1(new_n294), .C2(new_n293), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n224), .B1(new_n255), .B2(new_n256), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n460), .C1(new_n572), .C2(KEYINPUT4), .ZN(new_n573));
  OAI21_X1  g0373(.A(G250), .B1(new_n293), .B2(new_n294), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n258), .B1(new_n574), .B2(KEYINPUT4), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n262), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n476), .A2(G257), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(new_n253), .A3(new_n475), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  INV_X1    g0379(.A(G107), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n212), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G97), .A2(G107), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n520), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT77), .A2(G97), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(KEYINPUT6), .A3(new_n580), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n292), .A2(new_n296), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n290), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n456), .A2(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n314), .A2(new_n212), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n578), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n213), .B(new_n262), .C1(new_n474), .C2(new_n472), .ZN(new_n599));
  OAI21_X1  g0399(.A(G244), .B1(new_n293), .B2(new_n294), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n569), .B1(G33), .B2(G283), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n569), .B1(new_n257), .B2(G250), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n571), .C1(new_n258), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n603), .B2(new_n262), .ZN(new_n604));
  AOI21_X1  g0404(.A(G169), .B1(new_n604), .B2(new_n475), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n576), .A2(new_n475), .A3(new_n577), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n607), .A2(KEYINPUT79), .A3(G200), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT79), .B1(new_n607), .B2(G200), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n591), .A2(new_n597), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n604), .A2(G190), .A3(new_n475), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n606), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n513), .A2(new_n565), .A3(new_n568), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n454), .A2(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n545), .A2(new_n558), .ZN(new_n617));
  OR3_X1    g0417(.A1(new_n503), .A2(new_n560), .A3(new_n563), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n614), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT83), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n512), .A2(new_n503), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n483), .A3(new_n484), .A4(new_n481), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT83), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n565), .A2(new_n624), .A3(new_n614), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n545), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n545), .A2(new_n606), .A3(new_n558), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n545), .A2(new_n606), .A3(new_n558), .A4(KEYINPUT26), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n453), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n321), .A2(new_n325), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n425), .A2(new_n426), .B1(new_n415), .B2(new_n447), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n343), .A2(new_n344), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n374), .A2(new_n377), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n363), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n642), .B(KEYINPUT84), .Z(G369));
  INV_X1    g0443(.A(G13), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n203), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT27), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(G213), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n622), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n564), .B1(new_n503), .B2(new_n653), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n503), .B2(new_n512), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(new_n654), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n466), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n485), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n485), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n568), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n653), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n485), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n654), .B1(new_n658), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT86), .Z(G399));
  INV_X1    g0470(.A(new_n207), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G1), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n461), .A2(new_n215), .A3(new_n518), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n235), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n633), .A2(new_n666), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n565), .A2(new_n623), .A3(new_n614), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n632), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(new_n666), .ZN(new_n684));
  AOI211_X1 g0484(.A(KEYINPUT87), .B(new_n653), .C1(new_n632), .C2(new_n682), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n680), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT31), .B1(new_n615), .B2(new_n653), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n542), .A2(new_n561), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n482), .A4(new_n604), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n482), .A2(new_n604), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n542), .A2(new_n561), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n542), .A2(new_n566), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n253), .A3(new_n511), .A4(new_n607), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n653), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(G330), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n687), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n677), .B1(new_n704), .B2(G1), .ZN(G364));
  NAND2_X1  g0505(.A1(new_n662), .A2(new_n663), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT88), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n674), .B1(G45), .B2(new_n645), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n665), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n231), .B1(G20), .B2(new_n286), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n204), .A2(new_n253), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(G190), .A3(new_n562), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n226), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n253), .A2(new_n562), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n338), .A2(G20), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G159), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n295), .B(new_n715), .C1(KEYINPUT32), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n712), .A2(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n338), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n723), .B1(KEYINPUT32), .B2(new_n722), .C1(new_n221), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n562), .A2(G179), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(G20), .A3(G190), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n210), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n717), .A2(G190), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n204), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n719), .A2(new_n728), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n733), .A2(G97), .B1(G107), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n713), .A2(new_n338), .A3(new_n562), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n223), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n724), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n233), .ZN(new_n742));
  NOR4_X1   g0542(.A1(new_n727), .A2(new_n730), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n737), .A2(G311), .B1(G329), .B2(new_n721), .ZN(new_n744));
  INV_X1    g0544(.A(new_n714), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G322), .ZN(new_n746));
  INV_X1    g0546(.A(G294), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n744), .B(new_n746), .C1(new_n747), .C2(new_n732), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n729), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n725), .A2(G326), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT33), .B(G317), .Z(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n295), .B1(new_n741), .B2(new_n752), .C1(new_n734), .C2(new_n753), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n711), .B1(new_n743), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT89), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n709), .B1(new_n662), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n711), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n671), .A2(new_n257), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G45), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(new_n236), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n248), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G116), .B2(new_n207), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n671), .A2(new_n295), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G355), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n756), .B(new_n762), .C1(new_n764), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n710), .A2(new_n773), .ZN(G396));
  INV_X1    g0574(.A(new_n447), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n653), .A2(new_n437), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n451), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n678), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n778), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n633), .A2(new_n666), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n703), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT95), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n708), .B1(new_n782), .B2(new_n703), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n711), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n745), .A2(G143), .B1(G150), .B2(new_n740), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n789), .B2(new_n726), .C1(new_n301), .C2(new_n738), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT34), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n734), .A2(new_n233), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n295), .B1(new_n721), .B2(G132), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(KEYINPUT94), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n221), .B2(new_n729), .C1(new_n226), .C2(new_n732), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n737), .A2(G116), .B1(G283), .B2(new_n740), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n295), .B1(new_n799), .B2(KEYINPUT93), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n745), .A2(G294), .B1(G311), .B2(new_n721), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n801), .B1(new_n210), .B2(new_n734), .C1(new_n212), .C2(new_n732), .ZN(new_n802));
  INV_X1    g0602(.A(new_n729), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n800), .B(new_n802), .C1(G107), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT93), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n805), .B2(new_n798), .C1(new_n749), .C2(new_n726), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n787), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n780), .A2(new_n758), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n807), .A2(new_n709), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n711), .A2(new_n757), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(G77), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n786), .A2(new_n812), .ZN(G384));
  INV_X1    g0613(.A(KEYINPUT39), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n341), .A2(KEYINPUT98), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n323), .A2(new_n651), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n287), .B2(new_n320), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT98), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(new_n323), .C1(new_n337), .C2(new_n340), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT99), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n817), .A2(new_n823), .A3(new_n341), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT99), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT37), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n635), .A2(new_n638), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n816), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT38), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n651), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n309), .B1(KEYINPUT16), .B2(new_n308), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n319), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n327), .C2(new_n345), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n287), .B2(new_n831), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n341), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n824), .B1(new_n836), .B2(new_n823), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n814), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n427), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n425), .A2(KEYINPUT97), .A3(new_n426), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n653), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n834), .A2(new_n837), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n837), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n839), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n426), .A2(new_n653), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(new_n415), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n419), .A2(new_n427), .ZN(new_n854));
  INV_X1    g0654(.A(new_n852), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n843), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n775), .A2(new_n653), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n781), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n851), .A2(new_n859), .B1(new_n635), .B2(new_n651), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n680), .B(new_n453), .C1(new_n686), .C2(new_n679), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n641), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n861), .B(new_n863), .Z(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n834), .B2(new_n837), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n838), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT100), .B1(new_n698), .B2(new_n701), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n697), .A2(new_n869), .A3(KEYINPUT31), .A4(new_n653), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n688), .B2(new_n698), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n843), .A2(new_n853), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n854), .A2(new_n855), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n876), .A3(new_n780), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n865), .B1(new_n867), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n856), .A2(new_n872), .A3(new_n778), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT40), .B(new_n879), .C1(new_n830), .C2(new_n838), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n880), .A3(G330), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n872), .A2(new_n663), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n454), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n878), .A2(new_n880), .A3(new_n873), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n454), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n864), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n203), .B2(new_n645), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n215), .B1(new_n587), .B2(KEYINPUT35), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n232), .C1(KEYINPUT35), .C2(new_n587), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n235), .A2(new_n223), .A3(new_n299), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT96), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(G50), .B2(new_n233), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n644), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n891), .A3(new_n895), .ZN(G367));
  NOR2_X1   g0696(.A1(new_n244), .A2(new_n766), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n763), .B1(new_n207), .B2(new_n432), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n738), .A2(new_n221), .B1(new_n789), .B2(new_n720), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n295), .B(new_n899), .C1(G159), .C2(new_n740), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n735), .A2(G77), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n803), .A2(G58), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n745), .A2(G150), .B1(G143), .B2(new_n725), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n233), .B2(new_n732), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n732), .A2(new_n580), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n737), .A2(G283), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n721), .A2(G317), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n725), .A2(G311), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n729), .A2(new_n215), .ZN(new_n913));
  AOI22_X1  g0713(.A1(KEYINPUT46), .A2(new_n913), .B1(new_n740), .B2(G294), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n734), .A2(new_n461), .B1(KEYINPUT46), .B2(new_n913), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n915), .A2(new_n257), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n469), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n714), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n907), .A2(new_n908), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT47), .Z(new_n921));
  OAI221_X1 g0721(.A(new_n708), .B1(new_n897), .B2(new_n898), .C1(new_n921), .C2(new_n787), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  INV_X1    g0723(.A(new_n550), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n653), .B1(new_n924), .B2(new_n555), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n617), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n545), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n923), .B1(new_n760), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n645), .A2(G45), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G1), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n668), .B(new_n657), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n704), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n657), .A2(new_n667), .ZN(new_n933));
  INV_X1    g0733(.A(new_n654), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n614), .B1(new_n611), .B2(new_n666), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n606), .A2(new_n653), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT44), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n938), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT45), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n657), .A2(new_n665), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n704), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n672), .B(KEYINPUT41), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n930), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT42), .Z(new_n952));
  OAI22_X1  g0752(.A1(new_n936), .A2(new_n622), .B1(new_n605), .B2(new_n598), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n666), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n945), .A2(new_n938), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT101), .Z(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n955), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n928), .B1(new_n949), .B2(new_n960), .ZN(G387));
  NAND2_X1  g0761(.A1(new_n931), .A2(new_n930), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n738), .A2(new_n233), .B1(new_n221), .B2(new_n714), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n732), .A2(new_n432), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n720), .A2(new_n356), .B1(new_n734), .B2(new_n212), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n295), .B(new_n966), .C1(new_n429), .C2(new_n740), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n725), .A2(G159), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n803), .A2(G77), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n965), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n737), .A2(new_n469), .B1(G311), .B2(new_n740), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n745), .A2(G317), .ZN(new_n972));
  XNOR2_X1  g0772(.A(KEYINPUT105), .B(G322), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n971), .B(new_n972), .C1(new_n726), .C2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n753), .B2(new_n732), .C1(new_n747), .C2(new_n729), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT49), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n735), .A2(G116), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n721), .A2(G326), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n978), .A2(new_n295), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n976), .A2(new_n977), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n970), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n711), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n771), .A2(new_n675), .B1(new_n580), .B2(new_n671), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT104), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n313), .A2(KEYINPUT50), .A3(G50), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n675), .ZN(new_n988));
  NAND2_X1  g0788(.A1(G68), .A2(G77), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT50), .B1(new_n313), .B2(G50), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n988), .A2(new_n767), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n765), .B(new_n991), .C1(new_n241), .C2(new_n767), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n709), .B1(new_n993), .B2(new_n763), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n984), .B(new_n994), .C1(new_n658), .C2(new_n760), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n672), .B1(new_n704), .B2(new_n931), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n962), .B(new_n995), .C1(new_n932), .C2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT106), .Z(G393));
  NOR2_X1   g0798(.A1(new_n941), .A2(new_n943), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n945), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n672), .B(new_n946), .C1(new_n1000), .C2(new_n932), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n930), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n938), .A2(new_n760), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n745), .A2(G311), .B1(G317), .B2(new_n725), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n257), .B(new_n1005), .C1(G116), .C2(new_n733), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n747), .B2(new_n738), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n741), .A2(new_n918), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n729), .A2(new_n753), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n720), .A2(new_n973), .B1(new_n734), .B2(new_n580), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G143), .A2(new_n721), .B1(new_n735), .B2(G87), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n257), .C1(new_n233), .C2(new_n729), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(KEYINPUT107), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1013), .A2(KEYINPUT107), .B1(G77), .B2(new_n733), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n714), .A2(new_n301), .B1(new_n356), .B2(new_n726), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT51), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(new_n313), .C2(new_n738), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1014), .B(new_n1018), .C1(G50), .C2(new_n740), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n711), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n763), .B1(new_n207), .B2(new_n461), .C1(new_n251), .C2(new_n766), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n708), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT108), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1003), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1001), .A2(new_n1002), .A3(new_n1025), .ZN(G390));
  OAI211_X1 g0826(.A(G330), .B(new_n780), .C1(new_n700), .C2(new_n702), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n856), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n882), .A2(new_n780), .A3(new_n876), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(new_n781), .B2(new_n858), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1027), .A2(new_n856), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n780), .B1(new_n684), .B2(new_n685), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n858), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(KEYINPUT109), .A3(new_n858), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT110), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n874), .A2(new_n1038), .A3(new_n875), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n874), .B2(new_n875), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n883), .A2(new_n778), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1030), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT111), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n883), .B2(new_n454), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n882), .A2(new_n453), .A3(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n641), .A3(new_n862), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT112), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT37), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n825), .B1(new_n820), .B2(KEYINPUT37), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n824), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n829), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n846), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT39), .B1(new_n1054), .B2(new_n848), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n849), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1055), .A2(new_n1056), .B1(new_n844), .B2(new_n859), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1035), .A2(new_n1058), .A3(new_n1036), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n844), .B1(new_n1054), .B2(new_n848), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1027), .A2(new_n856), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1057), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1029), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n844), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n830), .B2(new_n838), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1032), .A2(KEYINPUT109), .A3(new_n858), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT109), .B1(new_n1032), .B2(new_n858), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1069), .B2(new_n1058), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n859), .A2(new_n844), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n839), .B2(new_n849), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1048), .A2(new_n1063), .A3(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1062), .B(new_n1041), .C1(new_n1068), .C2(new_n1067), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n781), .A2(new_n858), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n863), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1070), .A2(new_n1072), .A3(new_n1031), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1029), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1081), .B(KEYINPUT112), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1074), .A2(new_n1084), .A3(new_n672), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT113), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT113), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1074), .A2(new_n1084), .A3(new_n1087), .A4(new_n672), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1073), .A2(new_n1063), .A3(new_n930), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n757), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  AOI22_X1  g0892(.A1(new_n737), .A2(new_n1092), .B1(G128), .B2(new_n725), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n789), .B2(new_n741), .C1(new_n301), .C2(new_n732), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n295), .B1(new_n745), .B2(G132), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n221), .B2(new_n734), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n721), .A2(G125), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n729), .A2(new_n356), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n720), .A2(new_n747), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1102), .A2(new_n792), .A3(new_n730), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n295), .C1(new_n580), .C2(new_n741), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n732), .A2(new_n223), .B1(new_n714), .B2(new_n215), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n738), .A2(new_n461), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n726), .A2(new_n753), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n711), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n708), .B1(new_n429), .B2(new_n811), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT114), .Z(new_n1111));
  NAND3_X1  g0911(.A1(new_n1091), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1090), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1089), .A2(new_n1114), .ZN(G378));
  NAND2_X1  g0915(.A1(new_n831), .A2(new_n360), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n378), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n378), .A2(new_n1118), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1117), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n378), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT117), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n1119), .A3(new_n1116), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1123), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n881), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1129), .A2(new_n878), .A3(new_n880), .A4(G330), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n861), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n861), .A3(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n930), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1129), .A2(new_n757), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n810), .A2(new_n221), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n734), .A2(new_n226), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G283), .B2(new_n721), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n969), .C1(new_n212), .C2(new_n741), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n732), .A2(new_n233), .B1(new_n215), .B2(new_n726), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT116), .Z(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G107), .C2(new_n745), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n432), .B2(new_n738), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1147), .A2(G41), .A3(new_n257), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n221), .B1(new_n293), .B2(G41), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n733), .A2(G150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n745), .A2(G128), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n737), .A2(G137), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n725), .A2(G125), .B1(new_n803), .B2(new_n1092), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G132), .B2(new_n740), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT59), .ZN(new_n1157));
  AOI21_X1  g0957(.A(G33), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G41), .B1(new_n721), .B2(G124), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n301), .C2(new_n734), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n711), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1139), .A2(new_n708), .A3(new_n1140), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1138), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1073), .A2(new_n1063), .A3(new_n1079), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1136), .A2(new_n1135), .B1(new_n1167), .B2(new_n1080), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n672), .B1(new_n1168), .B2(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1167), .B2(new_n1080), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1135), .A2(KEYINPUT118), .A3(new_n1136), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT118), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1133), .A2(new_n1173), .A3(new_n1134), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1166), .B1(new_n1169), .B2(new_n1175), .ZN(G375));
  NAND2_X1  g0976(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1081), .A3(new_n948), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1058), .A2(new_n758), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n295), .B1(new_n738), .B2(new_n580), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n964), .B1(G283), .B2(new_n745), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT119), .Z(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n901), .C1(new_n749), .C2(new_n720), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(G97), .C2(new_n803), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n215), .B2(new_n741), .C1(new_n747), .C2(new_n726), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n737), .A2(G150), .B1(new_n740), .B2(new_n1092), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n221), .B2(new_n732), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1141), .B(new_n1187), .C1(G159), .C2(new_n803), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n725), .A2(G132), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n745), .A2(G137), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n295), .B1(new_n721), .B2(G128), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n787), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1179), .A2(new_n1193), .A3(new_n709), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n810), .A2(new_n233), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1079), .A2(new_n930), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1178), .A2(new_n1196), .ZN(G381));
  NAND2_X1  g0997(.A1(new_n1085), .A2(new_n1114), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1167), .A2(new_n1080), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1137), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n673), .B1(new_n1201), .B2(new_n1170), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1165), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1204), .B2(KEYINPUT120), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(KEYINPUT120), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G387), .A2(G390), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  OR2_X1    g1008(.A1(G381), .A2(G384), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(G407));
  INV_X1    g1011(.A(G213), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1206), .B2(new_n652), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G407), .ZN(G409));
  AND2_X1   g1014(.A1(G393), .A2(G396), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(new_n1208), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1216), .A2(KEYINPUT123), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(KEYINPUT123), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  INV_X1    g1020(.A(G390), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(G387), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n949), .A2(new_n960), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1223), .A2(KEYINPUT124), .A3(new_n928), .A4(G390), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(G387), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1216), .B1(G387), .B2(new_n1221), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1223), .A2(new_n928), .A3(G390), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1137), .A2(new_n1200), .A3(new_n948), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT121), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1168), .A2(KEYINPUT121), .A3(new_n948), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1172), .A2(new_n930), .A3(new_n1174), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1164), .A4(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G378), .A2(new_n1204), .B1(new_n1237), .B2(new_n1199), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1212), .A2(G343), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n673), .B1(new_n1177), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1081), .C1(new_n1241), .C2(new_n1177), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1196), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(G384), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT63), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT63), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1113), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G375), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT121), .B1(new_n1168), .B2(new_n948), .ZN(new_n1252));
  AND4_X1   g1052(.A1(KEYINPUT121), .A2(new_n1137), .A3(new_n1200), .A4(new_n948), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1236), .A2(new_n1164), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1198), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1249), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1239), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G378), .A2(new_n1204), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1237), .A2(new_n1199), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(KEYINPUT122), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1239), .A2(G2897), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1245), .B(new_n1263), .Z(new_n1264));
  AOI21_X1  g1064(.A(new_n1248), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1257), .A2(new_n1258), .A3(new_n1245), .A4(new_n1261), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1231), .B(new_n1247), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1219), .A2(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1270), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1245), .B(new_n1263), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1240), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1269), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1277), .ZN(G405));
  OAI21_X1  g1078(.A(new_n1259), .B1(new_n1204), .B2(new_n1198), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1245), .A2(KEYINPUT126), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1279), .B(new_n1280), .Z(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1269), .ZN(G402));
endmodule


