//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G127gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  AOI211_X1 g008(.A(KEYINPUT1), .B(G127gat), .C1(new_n203), .C2(new_n205), .ZN(new_n210));
  OAI21_X1  g009(.A(G134gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n207), .B(G127gat), .C1(new_n212), .C2(KEYINPUT1), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT76), .B1(new_n219), .B2(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT76), .ZN(new_n221));
  INV_X1    g020(.A(G141gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(G141gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  OR3_X1    g025(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n225), .A2(KEYINPUT77), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n220), .A2(new_n223), .A3(new_n229), .A4(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n224), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n219), .A2(G141gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n226), .B1(KEYINPUT75), .B2(KEYINPUT2), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n232), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n226), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n218), .B1(KEYINPUT3), .B2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n228), .A2(new_n230), .B1(new_n236), .B2(new_n240), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT78), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND4_X1   g045(.A1(KEYINPUT78), .A2(new_n231), .A3(new_n245), .A4(new_n241), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT4), .B1(new_n218), .B2(new_n244), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n248), .A2(new_n251), .A3(new_n255), .A4(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n211), .A3(new_n217), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n218), .A2(new_n244), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT5), .B1(new_n260), .B2(new_n252), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G1gat), .B(G29gat), .Z(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n253), .B2(KEYINPUT5), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(KEYINPUT81), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n268), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n261), .B1(new_n254), .B2(new_n256), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n273), .B2(new_n269), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(new_n275), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT6), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G29gat), .ZN(new_n282));
  INV_X1    g081(.A(G36gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT14), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT14), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G29gat), .B2(G36gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G29gat), .A2(G36gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT15), .ZN(new_n289));
  INV_X1    g088(.A(G43gat), .ZN(new_n290));
  INV_X1    g089(.A(G50gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G43gat), .A2(G50gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n296));
  NAND3_X1  g095(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n297));
  OR2_X1    g096(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n290), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n289), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n297), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n295), .B(new_n296), .C1(new_n303), .C2(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT93), .ZN(new_n305));
  INV_X1    g104(.A(G22gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G15gat), .ZN(new_n307));
  INV_X1    g106(.A(G15gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G22gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT16), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G1gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G8gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(KEYINPUT94), .ZN(new_n316));
  AND4_X1   g115(.A1(KEYINPUT94), .A2(new_n307), .A3(new_n309), .A4(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT94), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G8gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n315), .A2(KEYINPUT94), .A3(new_n314), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n312), .A4(new_n311), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n302), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n294), .B1(new_n324), .B2(new_n288), .ZN(new_n325));
  INV_X1    g124(.A(new_n294), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n297), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT17), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n301), .B1(new_n331), .B2(new_n290), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n326), .B1(new_n332), .B2(new_n297), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT93), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n295), .A4(new_n296), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n305), .A2(new_n323), .A3(new_n328), .A4(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n318), .A3(new_n322), .A4(new_n295), .ZN(new_n337));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT18), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n337), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n338), .B(KEYINPUT13), .Z(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n337), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n336), .A2(KEYINPUT95), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT95), .B1(new_n336), .B2(new_n347), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n342), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G169gat), .B(G197gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT90), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(G113gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(new_n222), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n352), .B(new_n204), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n356), .A2(new_n359), .A3(KEYINPUT12), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT12), .B1(new_n356), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n350), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n336), .A2(new_n347), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n336), .A2(new_n347), .A3(KEYINPUT95), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n340), .A2(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G230gat), .A2(G233gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(G85gat), .A2(G92gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G99gat), .A2(G106gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT8), .ZN(new_n380));
  OR2_X1    g179(.A1(G85gat), .A2(G92gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n379), .ZN(new_n383));
  NOR2_X1   g182(.A1(G99gat), .A2(G106gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT98), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(G99gat), .A2(G106gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT98), .B1(new_n387), .B2(new_n379), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n378), .B(new_n382), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n380), .A2(new_n376), .A3(new_n381), .A4(new_n377), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n383), .B2(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(KEYINPUT98), .A3(new_n379), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT99), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n390), .A2(new_n395), .A3(new_n391), .A4(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT9), .ZN(new_n398));
  INV_X1    g197(.A(G71gat), .ZN(new_n399));
  INV_X1    g198(.A(G78gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT96), .ZN(new_n402));
  XOR2_X1   g201(.A(G57gat), .B(G64gat), .Z(new_n403));
  AOI21_X1  g202(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G71gat), .B(G78gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G64gat), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(G57gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(G57gat), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(new_n413), .B1(new_n404), .B2(new_n405), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n408), .A3(new_n402), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n407), .A2(new_n409), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n414), .B2(new_n402), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT102), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n390), .A2(KEYINPUT102), .A3(new_n391), .A4(new_n392), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n389), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT10), .B1(new_n417), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT10), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n416), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n397), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n373), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n389), .A2(new_n424), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n416), .B1(new_n433), .B2(new_n422), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n394), .A2(new_n396), .B1(new_n410), .B2(new_n415), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n434), .A2(new_n435), .A3(new_n373), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G120gat), .B(G148gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G176gat), .B(G204gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n432), .A2(KEYINPUT103), .A3(new_n437), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n432), .B2(new_n437), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G155gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G183gat), .B(G211gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G231gat), .ZN(new_n453));
  INV_X1    g252(.A(G233gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n420), .B2(KEYINPUT21), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT21), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n416), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n214), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n416), .B2(new_n457), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT21), .B(new_n455), .C1(new_n410), .C2(new_n415), .ZN(new_n462));
  OAI21_X1  g261(.A(G127gat), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n420), .A2(KEYINPUT21), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n323), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n460), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n452), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n460), .A2(new_n463), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n464), .A2(new_n323), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(new_n452), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n335), .A2(new_n328), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n397), .A2(KEYINPUT100), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT100), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n394), .A2(new_n478), .A3(new_n396), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n305), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n325), .A2(new_n327), .ZN(new_n481));
  AND2_X1   g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n397), .A2(new_n481), .B1(KEYINPUT41), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G134gat), .B(G162gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n482), .A2(KEYINPUT41), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT97), .Z(new_n489));
  XOR2_X1   g288(.A(G190gat), .B(G218gat), .Z(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT101), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n489), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n485), .B1(new_n480), .B2(new_n483), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n483), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n484), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n497), .B2(new_n486), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n475), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n448), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n274), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n263), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT6), .A4(new_n272), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n280), .A2(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G211gat), .B(G218gat), .Z(new_n507));
  INV_X1    g306(.A(KEYINPUT22), .ZN(new_n508));
  NAND2_X1  g307(.A1(G211gat), .A2(G218gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n507), .A2(KEYINPUT71), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT70), .B(G197gat), .ZN(new_n511));
  INV_X1    g310(.A(G204gat), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n510), .A3(new_n513), .A4(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G226gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n454), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(KEYINPUT29), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G169gat), .ZN(new_n526));
  INV_X1    g325(.A(G176gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n526), .A2(new_n527), .B1(new_n529), .B2(KEYINPUT23), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n528), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(G176gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G183gat), .ZN(new_n538));
  INV_X1    g337(.A(G190gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT67), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(KEYINPUT67), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT25), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n538), .A2(new_n539), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G183gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n539), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(KEYINPUT28), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT26), .B1(new_n528), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(new_n526), .A3(new_n527), .A4(KEYINPUT68), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n555), .C1(new_n526), .C2(new_n527), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n557), .A3(new_n539), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n540), .B(new_n541), .C1(new_n548), .C2(KEYINPUT24), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT65), .B(G169gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n535), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n533), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT72), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n547), .A2(new_n559), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n525), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n523), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n521), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n523), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n565), .A2(new_n524), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n520), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n520), .B1(new_n569), .B2(new_n571), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n521), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT37), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G8gat), .B(G36gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT73), .ZN(new_n582));
  XNOR2_X1  g381(.A(G64gat), .B(G92gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT38), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n572), .A2(new_n576), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n566), .A2(new_n568), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n524), .ZN(new_n590));
  INV_X1    g389(.A(new_n571), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n520), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n576), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n595));
  INV_X1    g394(.A(new_n584), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n573), .B1(new_n572), .B2(new_n576), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT87), .B1(new_n598), .B2(new_n584), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n599), .A3(new_n577), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n588), .B1(new_n600), .B2(KEYINPUT38), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n506), .A2(new_n601), .A3(new_n279), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n517), .A2(new_n603), .A3(new_n519), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT3), .B1(new_n604), .B2(KEYINPUT84), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT84), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n517), .A2(new_n606), .A3(new_n603), .A4(new_n519), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n244), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT78), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n242), .B2(KEYINPUT3), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n244), .A2(KEYINPUT78), .A3(new_n245), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n521), .B1(new_n612), .B2(new_n603), .ZN(new_n613));
  OAI211_X1 g412(.A(G228gat), .B(G233gat), .C1(new_n608), .C2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT83), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n517), .A2(new_n603), .A3(new_n519), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n615), .B(new_n242), .C1(new_n616), .C2(KEYINPUT3), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n618));
  OAI211_X1 g417(.A(KEYINPUT83), .B(new_n618), .C1(new_n604), .C2(new_n244), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n603), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n520), .ZN(new_n622));
  NAND2_X1  g421(.A1(G228gat), .A2(G233gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n614), .A2(new_n624), .A3(G22gat), .ZN(new_n625));
  AOI21_X1  g424(.A(G22gat), .B1(new_n614), .B2(new_n624), .ZN(new_n626));
  XNOR2_X1  g425(.A(G78gat), .B(G106gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n291), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n625), .A2(new_n626), .B1(KEYINPUT85), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n624), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n306), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n630), .B(KEYINPUT85), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n614), .A2(new_n624), .A3(G22gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n248), .A2(new_n251), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640));
  INV_X1    g439(.A(new_n252), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n268), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n258), .A2(new_n252), .A3(new_n259), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT39), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n639), .B2(new_n641), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT40), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n648), .A2(new_n649), .A3(new_n268), .A4(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT30), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n572), .A2(new_n652), .A3(new_n576), .A4(new_n584), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n596), .B1(new_n592), .B2(new_n593), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(KEYINPUT30), .A3(new_n587), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n651), .A2(new_n275), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n638), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n602), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n281), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n638), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n565), .A2(new_n218), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n565), .A2(new_n218), .ZN(new_n664));
  NAND2_X1  g463(.A1(G227gat), .A2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT64), .Z(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT32), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(G15gat), .B(G43gat), .Z(new_n671));
  XNOR2_X1  g470(.A(G71gat), .B(G99gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n667), .B(KEYINPUT32), .C1(new_n669), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n664), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n665), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n666), .A2(KEYINPUT34), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n679), .A2(KEYINPUT34), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n681), .A3(new_n676), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT36), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n658), .A2(new_n662), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n685), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n281), .A2(new_n659), .A3(new_n638), .A4(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT35), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n625), .A2(new_n626), .A3(new_n634), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n630), .A2(KEYINPUT85), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n633), .B2(new_n636), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT88), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n674), .A2(new_n681), .A3(new_n676), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n681), .B1(new_n674), .B2(new_n676), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n683), .A2(KEYINPUT88), .A3(new_n684), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n659), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n506), .A2(new_n279), .ZN(new_n703));
  AOI22_X1  g502(.A1(KEYINPUT35), .A2(new_n690), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n372), .B(new_n500), .C1(new_n688), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT104), .ZN(new_n706));
  INV_X1    g505(.A(new_n372), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n690), .A2(KEYINPUT35), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n658), .A2(new_n662), .A3(new_n687), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n500), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n281), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n312), .ZN(G1324gat));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n714), .ZN(new_n717));
  INV_X1    g516(.A(new_n659), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n314), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT16), .B(G8gat), .ZN(new_n720));
  AOI211_X1 g519(.A(new_n659), .B(new_n720), .C1(new_n706), .C2(new_n714), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT42), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n718), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n720), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(G1325gat));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n700), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n717), .A2(new_n308), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n687), .B1(new_n706), .B2(new_n714), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n308), .ZN(G1326gat));
  NAND2_X1  g530(.A1(new_n717), .A2(new_n661), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  NOR2_X1   g533(.A1(new_n495), .A2(new_n498), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(new_n448), .A3(new_n475), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n712), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(new_n282), .A3(new_n280), .A4(new_n279), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n688), .B2(new_n704), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n448), .B(KEYINPUT106), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n369), .A2(new_n370), .A3(new_n362), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n364), .A2(KEYINPUT105), .A3(new_n371), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n744), .A2(new_n475), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n660), .A2(new_n752), .A3(new_n661), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n718), .B1(new_n279), .B2(new_n280), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT107), .B1(new_n754), .B2(new_n638), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n753), .A2(new_n658), .A3(new_n755), .A4(new_n687), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n736), .B1(new_n756), .B2(new_n710), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n742), .B(new_n751), .C1(new_n757), .C2(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g557(.A(G29gat), .B1(new_n758), .B2(new_n281), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n759), .ZN(G1328gat));
  NAND3_X1  g559(.A1(new_n738), .A2(new_n283), .A3(new_n718), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n758), .B2(new_n659), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G36gat), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n758), .A2(new_n764), .A3(new_n659), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n762), .B(new_n763), .C1(new_n766), .C2(new_n767), .ZN(G1329gat));
  OAI21_X1  g567(.A(G43gat), .B1(new_n758), .B2(new_n687), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n738), .A2(new_n290), .A3(new_n728), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1330gat));
  OAI22_X1  g574(.A1(new_n758), .A2(new_n638), .B1(new_n330), .B2(new_n329), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n738), .A2(new_n661), .A3(new_n331), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT48), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n750), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n743), .A2(new_n499), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n756), .B2(new_n710), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n281), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT109), .B(G57gat), .Z(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n787), .A2(new_n659), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(G1333gat));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n687), .A2(new_n399), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n786), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n399), .B1(new_n787), .B2(new_n727), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(new_n799), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT110), .B1(new_n786), .B2(new_n797), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n801), .B(new_n796), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n802), .A2(new_n806), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n786), .A2(new_n661), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g608(.A(new_n446), .B1(new_n443), .B2(new_n444), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n783), .A2(new_n475), .A3(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n742), .B(new_n811), .C1(new_n757), .C2(KEYINPUT44), .ZN(new_n812));
  OAI21_X1  g611(.A(G85gat), .B1(new_n812), .B2(new_n281), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n756), .A2(new_n710), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n783), .A2(new_n475), .ZN(new_n815));
  AND4_X1   g614(.A1(KEYINPUT51), .A2(new_n814), .A3(new_n735), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT51), .B1(new_n757), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n281), .A2(G85gat), .A3(new_n810), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(G1336gat));
  NOR2_X1   g619(.A1(new_n659), .A2(G92gat), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n744), .B(new_n821), .C1(new_n816), .C2(new_n817), .ZN(new_n822));
  OAI21_X1  g621(.A(G92gat), .B1(new_n812), .B2(new_n659), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1337gat));
  OAI21_X1  g627(.A(G99gat), .B1(new_n812), .B2(new_n687), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n727), .A2(G99gat), .A3(new_n810), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n818), .B2(new_n830), .ZN(G1338gat));
  NOR2_X1   g630(.A1(new_n638), .A2(G106gat), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n744), .B(new_n832), .C1(new_n816), .C2(new_n817), .ZN(new_n833));
  OAI21_X1  g632(.A(G106gat), .B1(new_n812), .B2(new_n638), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1339gat));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n500), .A2(new_n840), .A3(new_n750), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n500), .B2(new_n750), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n373), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n430), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n427), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n430), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT55), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n373), .C1(new_n427), .C2(new_n431), .ZN(new_n851));
  INV_X1    g650(.A(new_n440), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT113), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n373), .B1(new_n429), .B2(new_n397), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n850), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n432), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n852), .A4(new_n851), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n851), .B(new_n852), .C1(new_n846), .C2(new_n848), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n855), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n445), .A2(new_n854), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n356), .A2(new_n359), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n338), .B1(new_n336), .B2(new_n337), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n344), .A2(new_n345), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n371), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n863), .A2(new_n736), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n868), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n448), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n750), .B2(new_n863), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(new_n736), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n843), .B1(new_n873), .B2(new_n475), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n280), .A2(new_n874), .A3(new_n279), .A4(new_n638), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n689), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n718), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n750), .A2(G113gat), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT114), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n659), .A3(new_n728), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n707), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1340gat));
  NAND2_X1  g682(.A1(new_n448), .A2(new_n202), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT115), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G120gat), .B1(new_n881), .B2(new_n743), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1341gat));
  INV_X1    g687(.A(new_n475), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n881), .A2(new_n214), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n876), .A2(new_n718), .A3(new_n889), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT116), .ZN(new_n892));
  AOI21_X1  g691(.A(G127gat), .B1(new_n891), .B2(KEYINPUT116), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1342gat));
  OAI21_X1  g693(.A(G134gat), .B1(new_n881), .B2(new_n736), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT69), .B(G134gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n659), .A2(new_n735), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n876), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n899), .B2(new_n896), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n876), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n898), .ZN(new_n902));
  OAI221_X1 g701(.A(new_n895), .B1(new_n896), .B2(new_n899), .C1(new_n901), .C2(new_n902), .ZN(G1343gat));
  AND2_X1   g702(.A1(new_n874), .A2(new_n661), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n686), .A2(new_n281), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n906), .A2(G141gat), .A3(new_n718), .A4(new_n707), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n686), .A2(new_n281), .A3(new_n718), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n638), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n863), .A2(new_n736), .A3(new_n868), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n364), .A2(new_n371), .B1(new_n861), .B2(new_n855), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(new_n445), .A3(new_n854), .A4(new_n860), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n735), .B1(new_n915), .B2(new_n871), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n916), .B2(KEYINPUT118), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n445), .A2(new_n854), .A3(new_n860), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n862), .B1(new_n746), .B2(new_n747), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n918), .A2(new_n919), .B1(new_n810), .B2(new_n868), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n920), .A2(KEYINPUT118), .A3(new_n736), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n889), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n912), .B1(new_n922), .B2(new_n843), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n874), .B2(new_n661), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G141gat), .B1(new_n925), .B2(new_n707), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT119), .B(new_n909), .C1(new_n923), .C2(new_n924), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n783), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n907), .B1(new_n931), .B2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G1344gat));
  NAND4_X1  g733(.A1(new_n904), .A2(new_n219), .A3(new_n448), .A4(new_n909), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n929), .A2(new_n448), .A3(new_n930), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n219), .A2(KEYINPUT59), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n909), .A2(new_n448), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n872), .A2(new_n736), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n475), .B1(new_n941), .B2(new_n913), .ZN(new_n942));
  INV_X1    g741(.A(new_n842), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n500), .A2(new_n840), .A3(new_n750), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n911), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n920), .A2(new_n736), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n475), .B1(new_n947), .B2(new_n913), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n448), .A2(new_n499), .A3(new_n372), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n661), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n946), .A2(KEYINPUT120), .B1(new_n950), .B2(new_n910), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n874), .A2(new_n952), .A3(new_n911), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n940), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n219), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n946), .A2(KEYINPUT120), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n950), .A2(new_n910), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n957), .A2(new_n953), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT121), .B1(new_n959), .B2(new_n940), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n939), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n935), .B1(new_n938), .B2(new_n961), .ZN(G1345gat));
  NAND2_X1  g761(.A1(new_n929), .A2(new_n930), .ZN(new_n963));
  OAI21_X1  g762(.A(G155gat), .B1(new_n963), .B2(new_n889), .ZN(new_n964));
  OR4_X1    g763(.A1(G155gat), .A2(new_n906), .A3(new_n718), .A4(new_n889), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1346gat));
  OAI21_X1  g765(.A(G162gat), .B1(new_n963), .B2(new_n736), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n718), .A2(G162gat), .A3(new_n736), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n906), .B2(new_n968), .ZN(G1347gat));
  AND2_X1   g768(.A1(new_n874), .A2(new_n281), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n661), .A2(new_n659), .A3(new_n685), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n562), .A3(new_n783), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n874), .A2(new_n638), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n659), .B1(new_n279), .B2(new_n280), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(new_n728), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G169gat), .B1(new_n977), .B2(new_n707), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT122), .ZN(G1348gat));
  NOR3_X1   g779(.A1(new_n977), .A2(new_n527), .A3(new_n743), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n972), .A2(new_n448), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n527), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(KEYINPUT123), .A3(new_n527), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(G1349gat));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n549), .A3(new_n475), .ZN(new_n988));
  OAI21_X1  g787(.A(G183gat), .B1(new_n977), .B2(new_n889), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n988), .A2(new_n989), .A3(KEYINPUT124), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n539), .A3(new_n735), .ZN(new_n992));
  OAI21_X1  g791(.A(G190gat), .B1(new_n977), .B2(new_n736), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n993), .A2(KEYINPUT61), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(KEYINPUT61), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1351gat));
  NAND2_X1  g795(.A1(new_n687), .A2(new_n975), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n997), .B1(new_n951), .B2(new_n953), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(G197gat), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n999), .A2(new_n1000), .A3(new_n707), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n686), .A2(new_n659), .A3(new_n638), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n970), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(new_n783), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1001), .B1(new_n1006), .B2(new_n1000), .ZN(G1352gat));
  AND3_X1   g806(.A1(new_n1003), .A2(new_n512), .A3(new_n448), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  OAI21_X1  g808(.A(G204gat), .B1(new_n999), .B2(new_n743), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1353gat));
  INV_X1    g810(.A(G211gat), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1005), .A2(new_n1012), .A3(new_n475), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n475), .ZN(new_n1014));
  AND4_X1   g813(.A1(KEYINPUT126), .A2(new_n1014), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  AOI22_X1  g816(.A1(new_n1014), .A2(new_n1017), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1013), .B1(new_n1015), .B2(new_n1018), .ZN(G1354gat));
  AND2_X1   g818(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n735), .B1(new_n998), .B2(KEYINPUT127), .ZN(new_n1021));
  OAI21_X1  g820(.A(G218gat), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g821(.A(G218gat), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1005), .A2(new_n1023), .A3(new_n735), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1022), .A2(new_n1024), .ZN(G1355gat));
endmodule


