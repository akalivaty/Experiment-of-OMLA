

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736;

  INV_X2 U374 ( .A(G953), .ZN(n724) );
  NOR2_X1 U375 ( .A1(n702), .A2(G902), .ZN(n453) );
  NOR2_X2 U376 ( .A1(G902), .A2(n705), .ZN(n500) );
  XNOR2_X2 U377 ( .A(n499), .B(n498), .ZN(n705) );
  NAND2_X2 U378 ( .A1(n389), .A2(n390), .ZN(n688) );
  AND2_X2 U379 ( .A1(n393), .A2(n394), .ZN(n389) );
  NAND2_X1 U380 ( .A1(n716), .A2(n723), .ZN(n696) );
  NOR2_X2 U381 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X2 U382 ( .A1(n602), .A2(n576), .ZN(n579) );
  XNOR2_X2 U383 ( .A(G478), .B(n500), .ZN(n540) );
  XOR2_X2 U384 ( .A(KEYINPUT38), .B(n559), .Z(n673) );
  XNOR2_X1 U385 ( .A(n696), .B(KEYINPUT2), .ZN(n425) );
  INV_X2 U386 ( .A(n657), .ZN(n580) );
  INV_X1 U387 ( .A(G125), .ZN(n382) );
  AND2_X2 U388 ( .A1(n425), .A2(n512), .ZN(n707) );
  NOR2_X1 U389 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U390 ( .A(n361), .B(KEYINPUT80), .ZN(n611) );
  AND2_X1 U391 ( .A1(n368), .A2(n367), .ZN(n553) );
  AND2_X1 U392 ( .A1(n732), .A2(n608), .ZN(n595) );
  AND2_X1 U393 ( .A1(n584), .A2(n583), .ZN(n637) );
  NOR2_X1 U394 ( .A1(n600), .A2(n587), .ZN(n588) );
  XNOR2_X1 U395 ( .A(n415), .B(KEYINPUT31), .ZN(n650) );
  OR2_X1 U396 ( .A1(n688), .A2(n384), .ZN(n383) );
  BUF_X1 U397 ( .A(n524), .Z(n559) );
  XNOR2_X1 U398 ( .A(n710), .B(n407), .ZN(n624) );
  XNOR2_X1 U399 ( .A(n506), .B(KEYINPUT16), .ZN(n412) );
  XNOR2_X1 U400 ( .A(n508), .B(n381), .ZN(n476) );
  XNOR2_X1 U401 ( .A(n352), .B(n441), .ZN(n503) );
  XNOR2_X1 U402 ( .A(n382), .B(G146), .ZN(n508) );
  INV_X2 U403 ( .A(G113), .ZN(n380) );
  INV_X2 U404 ( .A(G122), .ZN(n402) );
  NOR2_X1 U405 ( .A1(n667), .A2(n602), .ZN(n415) );
  XOR2_X1 U406 ( .A(KEYINPUT101), .B(n523), .Z(n676) );
  XNOR2_X1 U407 ( .A(G137), .B(G140), .ZN(n454) );
  XNOR2_X1 U408 ( .A(n442), .B(n429), .ZN(n428) );
  XNOR2_X1 U409 ( .A(n440), .B(G146), .ZN(n429) );
  XNOR2_X1 U410 ( .A(n503), .B(n432), .ZN(n442) );
  XNOR2_X1 U411 ( .A(n408), .B(n510), .ZN(n407) );
  XNOR2_X1 U412 ( .A(n509), .B(n409), .ZN(n408) );
  NAND2_X1 U413 ( .A1(n524), .A2(n672), .ZN(n522) );
  XNOR2_X1 U414 ( .A(n414), .B(KEYINPUT92), .ZN(n605) );
  XNOR2_X1 U415 ( .A(n476), .B(n377), .ZN(n479) );
  XNOR2_X1 U416 ( .A(n505), .B(n378), .ZN(n377) );
  XNOR2_X1 U417 ( .A(n379), .B(G143), .ZN(n378) );
  INV_X1 U418 ( .A(G122), .ZN(n379) );
  INV_X1 U419 ( .A(G134), .ZN(n435) );
  INV_X1 U420 ( .A(KEYINPUT28), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n522), .B(n355), .ZN(n573) );
  XNOR2_X1 U422 ( .A(n474), .B(G472), .ZN(n427) );
  BUF_X1 U423 ( .A(n527), .Z(n660) );
  XNOR2_X1 U424 ( .A(n406), .B(n357), .ZN(n405) );
  INV_X1 U425 ( .A(n503), .ZN(n413) );
  XNOR2_X1 U426 ( .A(n412), .B(n507), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n353), .ZN(n708) );
  XNOR2_X1 U428 ( .A(n457), .B(n722), .ZN(n365) );
  XNOR2_X1 U429 ( .A(G110), .B(G119), .ZN(n456) );
  NAND2_X1 U430 ( .A1(n707), .A2(G217), .ZN(n421) );
  XNOR2_X1 U431 ( .A(n398), .B(n356), .ZN(n397) );
  NAND2_X1 U432 ( .A1(n707), .A2(G475), .ZN(n398) );
  XNOR2_X1 U433 ( .A(n371), .B(KEYINPUT79), .ZN(n693) );
  NOR2_X1 U434 ( .A1(n736), .A2(n734), .ZN(n551) );
  XNOR2_X1 U435 ( .A(G140), .B(G131), .ZN(n480) );
  XNOR2_X1 U436 ( .A(G137), .B(G113), .ZN(n438) );
  XOR2_X1 U437 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n439) );
  INV_X1 U438 ( .A(KEYINPUT10), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n363), .B(n400), .ZN(n495) );
  NAND2_X1 U440 ( .A1(n724), .A2(G234), .ZN(n400) );
  XNOR2_X1 U441 ( .A(n399), .B(KEYINPUT69), .ZN(n363) );
  XNOR2_X1 U442 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n399) );
  XNOR2_X1 U443 ( .A(n511), .B(n410), .ZN(n409) );
  XNOR2_X1 U444 ( .A(n411), .B(KEYINPUT4), .ZN(n410) );
  INV_X1 U445 ( .A(KEYINPUT18), .ZN(n411) );
  OR2_X1 U446 ( .A1(n732), .A2(n608), .ZN(n609) );
  INV_X1 U447 ( .A(KEYINPUT102), .ZN(n372) );
  NOR2_X1 U448 ( .A1(n675), .A2(n575), .ZN(n373) );
  XNOR2_X1 U449 ( .A(n664), .B(n426), .ZN(n589) );
  INV_X1 U450 ( .A(KEYINPUT6), .ZN(n426) );
  AND2_X1 U451 ( .A1(n656), .A2(n564), .ZN(n565) );
  INV_X1 U452 ( .A(n655), .ZN(n564) );
  XNOR2_X1 U453 ( .A(G119), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U454 ( .A(n423), .B(n422), .ZN(n431) );
  XNOR2_X1 U455 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n422) );
  XNOR2_X1 U456 ( .A(n455), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U457 ( .A(G128), .B(KEYINPUT23), .ZN(n455) );
  XOR2_X1 U458 ( .A(KEYINPUT4), .B(G131), .Z(n437) );
  INV_X1 U459 ( .A(G146), .ZN(n450) );
  XNOR2_X1 U460 ( .A(n360), .B(n446), .ZN(n449) );
  XOR2_X1 U461 ( .A(G101), .B(G107), .Z(n446) );
  XNOR2_X1 U462 ( .A(n447), .B(n354), .ZN(n360) );
  OR2_X1 U463 ( .A1(n723), .A2(KEYINPUT2), .ZN(n371) );
  NAND2_X1 U464 ( .A1(n388), .A2(n591), .ZN(n384) );
  AND2_X1 U465 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U466 ( .A(n489), .B(n488), .ZN(n539) );
  NOR2_X1 U467 ( .A1(G902), .A2(n617), .ZN(n489) );
  XNOR2_X1 U468 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X1 U469 ( .A1(n542), .A2(n567), .ZN(n643) );
  NOR2_X1 U470 ( .A1(n539), .A2(n540), .ZN(n638) );
  INV_X1 U471 ( .A(n660), .ZN(n583) );
  XNOR2_X1 U472 ( .A(n403), .B(n358), .ZN(G57) );
  NAND2_X1 U473 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U474 ( .A1(n419), .A2(n404), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n419) );
  NAND2_X1 U476 ( .A1(n397), .A2(n404), .ZN(n396) );
  XNOR2_X1 U477 ( .A(n376), .B(n375), .ZN(n703) );
  XNOR2_X1 U478 ( .A(n702), .B(n701), .ZN(n375) );
  NAND2_X1 U479 ( .A1(n707), .A2(G469), .ZN(n376) );
  NOR2_X1 U480 ( .A1(n699), .A2(n700), .ZN(n366) );
  XOR2_X1 U481 ( .A(G101), .B(G116), .Z(n352) );
  XOR2_X1 U482 ( .A(n431), .B(n456), .Z(n353) );
  INV_X1 U483 ( .A(n602), .ZN(n388) );
  XOR2_X1 U484 ( .A(G110), .B(G104), .Z(n354) );
  XNOR2_X1 U485 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n355) );
  INV_X1 U486 ( .A(n591), .ZN(n395) );
  XOR2_X1 U487 ( .A(n619), .B(n618), .Z(n356) );
  XNOR2_X1 U488 ( .A(n472), .B(n445), .ZN(n357) );
  XOR2_X1 U489 ( .A(G902), .B(KEYINPUT15), .Z(n512) );
  NOR2_X1 U490 ( .A1(G952), .A2(n724), .ZN(n709) );
  INV_X1 U491 ( .A(n709), .ZN(n404) );
  XOR2_X1 U492 ( .A(n616), .B(KEYINPUT63), .Z(n358) );
  XOR2_X1 U493 ( .A(n620), .B(KEYINPUT67), .Z(n359) );
  NAND2_X1 U494 ( .A1(n650), .A2(n634), .ZN(n414) );
  XNOR2_X1 U495 ( .A(n428), .B(n721), .ZN(n472) );
  NAND2_X1 U496 ( .A1(n610), .A2(n609), .ZN(n361) );
  NAND2_X1 U497 ( .A1(n362), .A2(n436), .ZN(n490) );
  NAND2_X1 U498 ( .A1(n424), .A2(n435), .ZN(n362) );
  XNOR2_X1 U499 ( .A(n373), .B(n372), .ZN(n576) );
  NAND2_X1 U500 ( .A1(n374), .A2(n540), .ZN(n675) );
  XNOR2_X2 U501 ( .A(n364), .B(n413), .ZN(n710) );
  XNOR2_X1 U502 ( .A(n366), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U503 ( .A(n653), .ZN(n367) );
  NOR2_X1 U504 ( .A1(n538), .A2(n537), .ZN(n368) );
  NAND2_X1 U505 ( .A1(n369), .A2(n521), .ZN(n542) );
  XNOR2_X1 U506 ( .A(n520), .B(n370), .ZN(n369) );
  INV_X1 U507 ( .A(n539), .ZN(n374) );
  XNOR2_X2 U508 ( .A(n380), .B(G104), .ZN(n505) );
  NAND2_X1 U509 ( .A1(n385), .A2(n383), .ZN(n592) );
  NAND2_X1 U510 ( .A1(n602), .A2(n395), .ZN(n386) );
  NAND2_X1 U511 ( .A1(n688), .A2(n395), .ZN(n387) );
  NAND2_X1 U512 ( .A1(n391), .A2(n392), .ZN(n390) );
  NOR2_X1 U513 ( .A1(n658), .A2(n590), .ZN(n391) );
  INV_X1 U514 ( .A(n417), .ZN(n392) );
  NAND2_X1 U515 ( .A1(n658), .A2(n590), .ZN(n393) );
  NAND2_X1 U516 ( .A1(n417), .A2(n590), .ZN(n394) );
  XNOR2_X1 U517 ( .A(n396), .B(n359), .ZN(G60) );
  XNOR2_X2 U518 ( .A(n528), .B(KEYINPUT68), .ZN(n658) );
  XNOR2_X2 U519 ( .A(n453), .B(G469), .ZN(n529) );
  XNOR2_X1 U520 ( .A(n582), .B(KEYINPUT64), .ZN(n584) );
  AND2_X1 U521 ( .A1(n553), .A2(n552), .ZN(n554) );
  AND2_X2 U522 ( .A1(n566), .A2(n565), .ZN(n723) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(n527) );
  NAND2_X1 U524 ( .A1(n401), .A2(n585), .ZN(n600) );
  AND2_X1 U525 ( .A1(n401), .A2(n581), .ZN(n582) );
  XNOR2_X1 U526 ( .A(n579), .B(n578), .ZN(n401) );
  INV_X1 U527 ( .A(n573), .ZN(n567) );
  XNOR2_X2 U528 ( .A(n514), .B(n513), .ZN(n524) );
  XNOR2_X2 U529 ( .A(n402), .B(G107), .ZN(n504) );
  NAND2_X1 U530 ( .A1(n707), .A2(G472), .ZN(n406) );
  NOR2_X1 U531 ( .A1(n658), .A2(n416), .ZN(n601) );
  NAND2_X1 U532 ( .A1(n580), .A2(n664), .ZN(n416) );
  NAND2_X1 U533 ( .A1(n580), .A2(n589), .ZN(n417) );
  XNOR2_X1 U534 ( .A(n418), .B(KEYINPUT123), .ZN(G66) );
  INV_X1 U535 ( .A(n708), .ZN(n420) );
  INV_X1 U536 ( .A(n434), .ZN(n424) );
  XNOR2_X1 U537 ( .A(n434), .B(KEYINPUT17), .ZN(n509) );
  XNOR2_X2 U538 ( .A(n473), .B(n427), .ZN(n664) );
  XNOR2_X2 U539 ( .A(n490), .B(n437), .ZN(n721) );
  NOR2_X2 U540 ( .A1(n627), .A2(n709), .ZN(n629) );
  XNOR2_X1 U541 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X2 U542 ( .A(n594), .B(KEYINPUT35), .ZN(n732) );
  XOR2_X1 U543 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n430) );
  NAND2_X1 U544 ( .A1(n477), .A2(G210), .ZN(n432) );
  OR2_X1 U545 ( .A1(n597), .A2(n608), .ZN(n433) );
  XNOR2_X1 U546 ( .A(n460), .B(KEYINPUT25), .ZN(n461) );
  XNOR2_X1 U547 ( .A(n721), .B(n450), .ZN(n451) );
  INV_X1 U548 ( .A(KEYINPUT60), .ZN(n620) );
  XNOR2_X2 U549 ( .A(G128), .B(G143), .ZN(n434) );
  NAND2_X1 U550 ( .A1(n434), .A2(G134), .ZN(n436) );
  XNOR2_X1 U551 ( .A(n439), .B(n438), .ZN(n440) );
  NOR2_X1 U552 ( .A1(G953), .A2(G237), .ZN(n477) );
  XOR2_X1 U553 ( .A(KEYINPUT83), .B(KEYINPUT112), .Z(n444) );
  XNOR2_X1 U554 ( .A(KEYINPUT62), .B(KEYINPUT111), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U556 ( .A(n454), .ZN(n447) );
  NAND2_X1 U557 ( .A1(G227), .A2(n724), .ZN(n448) );
  XNOR2_X1 U558 ( .A(n449), .B(n448), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n452), .B(n451), .ZN(n702) );
  XNOR2_X2 U560 ( .A(n529), .B(KEYINPUT1), .ZN(n657) );
  XNOR2_X1 U561 ( .A(n476), .B(n454), .ZN(n722) );
  NAND2_X1 U562 ( .A1(G221), .A2(n495), .ZN(n457) );
  NOR2_X1 U563 ( .A1(n708), .A2(G902), .ZN(n462) );
  XOR2_X1 U564 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n459) );
  INV_X1 U565 ( .A(n512), .ZN(n615) );
  NAND2_X1 U566 ( .A1(G234), .A2(n615), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n459), .B(n458), .ZN(n468) );
  NAND2_X1 U568 ( .A1(n468), .A2(G217), .ZN(n460) );
  NAND2_X1 U569 ( .A1(G237), .A2(G234), .ZN(n463) );
  XNOR2_X1 U570 ( .A(n463), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U571 ( .A1(G952), .A2(n465), .ZN(n464) );
  XNOR2_X1 U572 ( .A(KEYINPUT86), .B(n464), .ZN(n686) );
  NOR2_X1 U573 ( .A1(G953), .A2(n686), .ZN(n568) );
  AND2_X1 U574 ( .A1(G902), .A2(n465), .ZN(n569) );
  NAND2_X1 U575 ( .A1(G953), .A2(n569), .ZN(n466) );
  NOR2_X1 U576 ( .A1(G900), .A2(n466), .ZN(n467) );
  NOR2_X1 U577 ( .A1(n568), .A2(n467), .ZN(n545) );
  NAND2_X1 U578 ( .A1(n468), .A2(G221), .ZN(n469) );
  XOR2_X1 U579 ( .A(KEYINPUT21), .B(n469), .Z(n661) );
  INV_X1 U580 ( .A(n661), .ZN(n575) );
  NOR2_X1 U581 ( .A1(n545), .A2(n575), .ZN(n470) );
  XNOR2_X1 U582 ( .A(n470), .B(KEYINPUT71), .ZN(n471) );
  NOR2_X1 U583 ( .A1(n527), .A2(n471), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT73), .B(KEYINPUT90), .ZN(n474) );
  NOR2_X1 U585 ( .A1(G902), .A2(n472), .ZN(n473) );
  NAND2_X1 U586 ( .A1(n518), .A2(n589), .ZN(n475) );
  XNOR2_X1 U587 ( .A(n475), .B(KEYINPUT105), .ZN(n501) );
  NAND2_X1 U588 ( .A1(n477), .A2(G214), .ZN(n478) );
  XNOR2_X1 U589 ( .A(n479), .B(n478), .ZN(n487) );
  XOR2_X1 U590 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n481) );
  XNOR2_X1 U591 ( .A(n481), .B(n480), .ZN(n485) );
  XOR2_X1 U592 ( .A(KEYINPUT12), .B(KEYINPUT93), .Z(n483) );
  XNOR2_X1 U593 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U594 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U595 ( .A(n485), .B(n484), .Z(n486) );
  XNOR2_X1 U596 ( .A(n487), .B(n486), .ZN(n617) );
  XNOR2_X1 U597 ( .A(KEYINPUT13), .B(G475), .ZN(n488) );
  XOR2_X1 U598 ( .A(KEYINPUT98), .B(n490), .Z(n492) );
  XNOR2_X1 U599 ( .A(n504), .B(G116), .ZN(n491) );
  XNOR2_X1 U600 ( .A(n492), .B(n491), .ZN(n499) );
  XOR2_X1 U601 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n494) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT99), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n497) );
  NAND2_X1 U604 ( .A1(G217), .A2(n495), .ZN(n496) );
  XOR2_X1 U605 ( .A(n497), .B(n496), .Z(n498) );
  NAND2_X1 U606 ( .A1(n539), .A2(n540), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT104), .B(n549), .Z(n644) );
  NAND2_X1 U608 ( .A1(n501), .A2(n644), .ZN(n502) );
  XNOR2_X1 U609 ( .A(KEYINPUT106), .B(n502), .ZN(n555) );
  XNOR2_X1 U610 ( .A(G110), .B(n504), .ZN(n507) );
  INV_X1 U611 ( .A(n505), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n508), .B(KEYINPUT85), .ZN(n510) );
  NAND2_X1 U613 ( .A1(G224), .A2(n724), .ZN(n511) );
  NOR2_X2 U614 ( .A1(n512), .A2(n624), .ZN(n514) );
  OR2_X1 U615 ( .A1(G902), .A2(G237), .ZN(n515) );
  NAND2_X1 U616 ( .A1(G210), .A2(n515), .ZN(n513) );
  NAND2_X1 U617 ( .A1(G214), .A2(n515), .ZN(n672) );
  NOR2_X1 U618 ( .A1(n555), .A2(n522), .ZN(n516) );
  XOR2_X1 U619 ( .A(KEYINPUT36), .B(n516), .Z(n517) );
  NOR2_X1 U620 ( .A1(n657), .A2(n517), .ZN(n653) );
  NAND2_X1 U621 ( .A1(n518), .A2(n664), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n519), .B(n430), .ZN(n520) );
  INV_X1 U623 ( .A(n529), .ZN(n521) );
  XOR2_X1 U624 ( .A(KEYINPUT100), .B(n638), .Z(n563) );
  NAND2_X1 U625 ( .A1(n549), .A2(n563), .ZN(n523) );
  NAND2_X1 U626 ( .A1(n643), .A2(n676), .ZN(n536) );
  NAND2_X1 U627 ( .A1(n536), .A2(KEYINPUT47), .ZN(n534) );
  NAND2_X1 U628 ( .A1(n664), .A2(n672), .ZN(n526) );
  XOR2_X1 U629 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n525) );
  XNOR2_X1 U630 ( .A(n526), .B(n525), .ZN(n530) );
  NAND2_X1 U631 ( .A1(n661), .A2(n527), .ZN(n528) );
  NOR2_X1 U632 ( .A1(n658), .A2(n529), .ZN(n604) );
  NAND2_X1 U633 ( .A1(n530), .A2(n604), .ZN(n546) );
  OR2_X1 U634 ( .A1(n545), .A2(n546), .ZN(n532) );
  INV_X1 U635 ( .A(n540), .ZN(n531) );
  NAND2_X1 U636 ( .A1(n539), .A2(n531), .ZN(n593) );
  NOR2_X1 U637 ( .A1(n532), .A2(n593), .ZN(n533) );
  NAND2_X1 U638 ( .A1(n559), .A2(n533), .ZN(n642) );
  NAND2_X1 U639 ( .A1(n534), .A2(n642), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n535), .B(KEYINPUT78), .ZN(n538) );
  NOR2_X1 U641 ( .A1(n536), .A2(KEYINPUT47), .ZN(n537) );
  NAND2_X1 U642 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U643 ( .A1(n677), .A2(n675), .ZN(n541) );
  XNOR2_X1 U644 ( .A(KEYINPUT41), .B(n541), .ZN(n687) );
  NOR2_X1 U645 ( .A1(n542), .A2(n687), .ZN(n543) );
  XNOR2_X1 U646 ( .A(KEYINPUT42), .B(n543), .ZN(n736) );
  INV_X1 U647 ( .A(n673), .ZN(n544) );
  OR2_X1 U648 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U649 ( .A(n548), .B(KEYINPUT39), .ZN(n562) );
  NOR2_X1 U650 ( .A1(n562), .A2(n549), .ZN(n550) );
  XNOR2_X1 U651 ( .A(KEYINPUT40), .B(n550), .ZN(n734) );
  XNOR2_X1 U652 ( .A(n551), .B(KEYINPUT46), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n554), .B(KEYINPUT48), .ZN(n566) );
  XOR2_X1 U654 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n558) );
  NOR2_X1 U655 ( .A1(n555), .A2(n580), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n556), .A2(n672), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n558), .B(n557), .ZN(n561) );
  INV_X1 U658 ( .A(n559), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n656) );
  NOR2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n655) );
  INV_X1 U661 ( .A(n568), .ZN(n571) );
  NOR2_X1 U662 ( .A1(G898), .A2(n724), .ZN(n712) );
  NAND2_X1 U663 ( .A1(n569), .A2(n712), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X2 U666 ( .A(n574), .B(KEYINPUT0), .ZN(n602) );
  XOR2_X1 U667 ( .A(KEYINPUT65), .B(KEYINPUT74), .Z(n577) );
  XNOR2_X1 U668 ( .A(KEYINPUT22), .B(n577), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n580), .A2(n664), .ZN(n581) );
  INV_X1 U670 ( .A(n589), .ZN(n585) );
  NOR2_X1 U671 ( .A1(n657), .A2(n660), .ZN(n586) );
  XNOR2_X1 U672 ( .A(n586), .B(KEYINPUT103), .ZN(n587) );
  XNOR2_X1 U673 ( .A(KEYINPUT32), .B(n588), .ZN(n733) );
  NOR2_X1 U674 ( .A1(n637), .A2(n733), .ZN(n597) );
  XOR2_X1 U675 ( .A(KEYINPUT82), .B(KEYINPUT33), .Z(n590) );
  XOR2_X1 U676 ( .A(KEYINPUT34), .B(KEYINPUT76), .Z(n591) );
  NOR2_X2 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n597), .A2(n595), .ZN(n596) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT72), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n598), .A2(n433), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n657), .A2(n660), .ZN(n599) );
  NOR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n630) );
  INV_X1 U684 ( .A(n630), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT91), .ZN(n667) );
  NOR2_X1 U686 ( .A1(n602), .A2(n664), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n634) );
  NAND2_X1 U688 ( .A1(n605), .A2(n676), .ZN(n606) );
  AND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n610) );
  NOR2_X2 U690 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U691 ( .A(KEYINPUT45), .ZN(n613) );
  XNOR2_X2 U692 ( .A(n614), .B(n613), .ZN(n716) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n695) );
  XNOR2_X1 U694 ( .A(KEYINPUT84), .B(KEYINPUT113), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT59), .B(KEYINPUT122), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n617), .B(KEYINPUT121), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n707), .A2(G210), .ZN(n626) );
  XOR2_X1 U698 ( .A(KEYINPUT55), .B(KEYINPUT81), .Z(n622) );
  XNOR2_X1 U699 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT56), .B(KEYINPUT120), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(G51) );
  XOR2_X1 U703 ( .A(G101), .B(n630), .Z(G3) );
  INV_X1 U704 ( .A(n644), .ZN(n646) );
  NOR2_X1 U705 ( .A1(n646), .A2(n634), .ZN(n631) );
  XOR2_X1 U706 ( .A(G104), .B(n631), .Z(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n633) );
  XNOR2_X1 U708 ( .A(G107), .B(KEYINPUT27), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(n636) );
  INV_X1 U710 ( .A(n638), .ZN(n651) );
  NOR2_X1 U711 ( .A1(n651), .A2(n634), .ZN(n635) );
  XOR2_X1 U712 ( .A(n636), .B(n635), .Z(G9) );
  XOR2_X1 U713 ( .A(n637), .B(G110), .Z(G12) );
  XOR2_X1 U714 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n640) );
  NAND2_X1 U715 ( .A1(n643), .A2(n638), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U717 ( .A(G128), .B(n641), .Z(G30) );
  XNOR2_X1 U718 ( .A(G143), .B(n642), .ZN(G45) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(G146), .ZN(G48) );
  NOR2_X1 U721 ( .A1(n646), .A2(n650), .ZN(n648) );
  XNOR2_X1 U722 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(G113), .B(n649), .ZN(G15) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(G116), .B(n652), .Z(G18) );
  XNOR2_X1 U727 ( .A(G125), .B(n653), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U729 ( .A(G134), .B(n655), .Z(G36) );
  XNOR2_X1 U730 ( .A(G140), .B(n656), .ZN(G42) );
  XOR2_X1 U731 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n670) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U739 ( .A(n670), .B(n669), .Z(n671) );
  NOR2_X1 U740 ( .A1(n687), .A2(n671), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n680) );
  INV_X1 U743 ( .A(n676), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n688), .A2(n681), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U752 ( .A1(n691), .A2(n724), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n716), .A2(KEYINPUT2), .ZN(n692) );
  XNOR2_X1 U754 ( .A(n694), .B(KEYINPUT77), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n701) );
  NOR2_X1 U758 ( .A1(n709), .A2(n703), .ZN(G54) );
  NAND2_X1 U759 ( .A1(G478), .A2(n707), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n709), .A2(n706), .ZN(G63) );
  XNOR2_X1 U762 ( .A(KEYINPUT125), .B(n710), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n720) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U766 ( .A1(n714), .A2(G898), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n715), .B(KEYINPUT124), .ZN(n718) );
  NAND2_X1 U768 ( .A1(n716), .A2(n724), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n727) );
  XOR2_X1 U772 ( .A(n727), .B(n723), .Z(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n726), .B(KEYINPUT126), .ZN(n731) );
  XNOR2_X1 U775 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n732), .B(G122), .ZN(G24) );
  XOR2_X1 U780 ( .A(n733), .B(G119), .Z(G21) );
  XNOR2_X1 U781 ( .A(G131), .B(KEYINPUT127), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(G33) );
  XOR2_X1 U783 ( .A(G137), .B(n736), .Z(G39) );
endmodule

