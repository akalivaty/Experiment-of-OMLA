//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(new_n203), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n213), .B1(new_n216), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  NAND2_X1  g0036(.A1(new_n201), .A2(G68), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n203), .A2(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G97), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G223), .A3(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G77), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n252), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT66), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n252), .A2(new_n253), .A3(new_n261), .A4(new_n257), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n247), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n264), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n270), .B2(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n263), .A2(G190), .A3(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n214), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT8), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G58), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(KEYINPUT67), .A3(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n208), .A3(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n279), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n208), .A3(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n201), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n279), .B1(G1), .B2(new_n208), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n201), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n276), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n295), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n287), .A2(new_n289), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n297), .B(KEYINPUT9), .C1(new_n298), .C2(new_n279), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n275), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n274), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n296), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n273), .A3(new_n303), .A4(new_n275), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n272), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n297), .B1(new_n298), .B2(new_n279), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n308), .C1(G179), .C2(new_n272), .ZN(new_n309));
  INV_X1    g0109(.A(new_n266), .ZN(new_n310));
  INV_X1    g0110(.A(G244), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n269), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n250), .A2(G238), .A3(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n250), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n316), .B2(new_n260), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G179), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n208), .A2(G33), .ZN(new_n321));
  OR3_X1    g0121(.A1(new_n320), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n281), .A2(new_n285), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT68), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n278), .ZN(new_n327));
  INV_X1    g0127(.A(new_n292), .ZN(new_n328));
  MUX2_X1   g0128(.A(new_n328), .B(new_n294), .S(G77), .Z(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n317), .A2(G169), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n319), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n327), .B(new_n329), .C1(new_n317), .C2(new_n335), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(KEYINPUT69), .B1(G190), .B2(new_n317), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND4_X1   g0139(.A1(new_n305), .A2(new_n309), .A3(new_n334), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n288), .A2(new_n341), .A3(G50), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n208), .B2(G68), .C1(new_n343), .C2(new_n321), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n341), .B1(new_n288), .B2(G50), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n278), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT11), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT12), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n203), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n328), .A2(new_n350), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n292), .A2(new_n348), .A3(new_n349), .A4(new_n203), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n292), .A2(new_n278), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n310), .B1(new_n269), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n361));
  OAI211_X1 g0161(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n268), .B1(new_n364), .B2(KEYINPUT70), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n362), .A3(new_n366), .A4(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n360), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n260), .A3(new_n367), .ZN(new_n372));
  INV_X1    g0172(.A(new_n360), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n368), .B2(new_n369), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  AOI211_X1 g0179(.A(KEYINPUT13), .B(new_n360), .C1(new_n365), .C2(new_n367), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(G169), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n380), .B2(new_n381), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n357), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G200), .B1(new_n380), .B2(new_n381), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n357), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n368), .B2(new_n369), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n370), .A2(new_n375), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n370), .A2(new_n375), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n251), .A2(G226), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n250), .B(new_n397), .C1(G223), .C2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n268), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n310), .B1(new_n269), .B2(new_n229), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n400), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n260), .ZN(new_n404));
  INV_X1    g0204(.A(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(G200), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n248), .A2(new_n208), .A3(new_n249), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n248), .A2(new_n410), .A3(new_n208), .A4(new_n249), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(G68), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(G58), .B(G68), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n279), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n412), .A2(new_n418), .A3(KEYINPUT16), .A4(new_n414), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT75), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n294), .A2(new_n286), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n292), .B2(new_n286), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n407), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n422), .A2(new_n424), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n404), .A2(new_n376), .A3(new_n405), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n306), .B1(new_n400), .B2(new_n401), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n422), .B2(new_n424), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT76), .B1(new_n439), .B2(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n429), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n340), .A2(new_n396), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n340), .A2(new_n396), .A3(new_n446), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G250), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n449));
  OAI211_X1 g0249(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n450));
  INV_X1    g0250(.A(G294), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n247), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n207), .A2(G45), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n260), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n452), .A2(new_n260), .B1(new_n456), .B2(G264), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n455), .A2(new_n268), .A3(G274), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n306), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G179), .B2(new_n459), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G116), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G20), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT23), .B1(new_n315), .B2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n315), .A2(KEYINPUT23), .A3(G20), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G87), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(KEYINPUT87), .B2(KEYINPUT22), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n250), .A2(new_n208), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT88), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n473));
  AOI21_X1  g0273(.A(G20), .B1(new_n248), .B2(new_n249), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT88), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n470), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n472), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT24), .ZN(new_n480));
  INV_X1    g0280(.A(new_n476), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n475), .B1(new_n474), .B2(new_n470), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n481), .A2(new_n482), .B1(KEYINPUT87), .B2(KEYINPUT22), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n468), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n279), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n207), .A2(G33), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n353), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT25), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n328), .B2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n315), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n493), .A2(G107), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n462), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n208), .C1(G33), .C2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT86), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G20), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n278), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n278), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(KEYINPUT20), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n328), .A2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n492), .B2(new_n504), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n455), .A2(new_n454), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n260), .A2(new_n265), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n456), .A2(G270), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G264), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n522));
  INV_X1    g0322(.A(G303), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n250), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n260), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n517), .A2(KEYINPUT21), .A3(G169), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n510), .B2(new_n511), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(G169), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n520), .A2(G179), .A3(new_n525), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n517), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n526), .A2(G200), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n520), .A2(G190), .A3(new_n525), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND4_X1   g0337(.A1(new_n527), .A2(new_n531), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n486), .B1(new_n485), .B2(new_n468), .ZN(new_n539));
  INV_X1    g0339(.A(new_n468), .ZN(new_n540));
  AOI211_X1 g0340(.A(KEYINPUT24), .B(new_n540), .C1(new_n483), .C2(new_n484), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n278), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n459), .A2(new_n335), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G190), .B2(new_n459), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n497), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT85), .B(G87), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n208), .B1(new_n363), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n208), .C1(new_n363), .C2(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n474), .A2(G68), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n321), .B2(new_n501), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n278), .B1(new_n292), .B2(new_n320), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n453), .A2(G250), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n260), .A2(new_n559), .B1(new_n265), .B2(new_n453), .ZN(new_n560));
  OAI211_X1 g0360(.A(G238), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n561));
  OAI211_X1 g0361(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n463), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(new_n260), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n493), .A2(G87), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  INV_X1    g0369(.A(new_n320), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n493), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n558), .A2(new_n571), .B1(new_n376), .B2(new_n564), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n306), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n567), .A2(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n499), .A2(new_n538), .A3(new_n545), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n579));
  XOR2_X1   g0379(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n250), .A2(KEYINPUT80), .A3(G250), .A4(G1698), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n500), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n260), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n455), .A2(new_n454), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(G257), .A3(new_n268), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n458), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT81), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n592), .A3(new_n458), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(new_n376), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n292), .A2(new_n501), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n492), .B2(new_n501), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n243), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n315), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(G20), .B1(G77), .B2(new_n288), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n409), .A2(G107), .A3(new_n411), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n605), .B2(new_n278), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n587), .A2(new_n591), .A3(new_n593), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n306), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n589), .A2(new_n592), .A3(new_n458), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n592), .B1(new_n589), .B2(new_n458), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT82), .A3(new_n376), .A4(new_n587), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n596), .A2(new_n607), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n606), .B1(new_n306), .B2(new_n608), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT83), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n613), .A4(new_n596), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n608), .A2(G200), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n606), .C1(new_n389), .C2(new_n608), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n575), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n448), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n386), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n395), .B2(new_n334), .ZN(new_n625));
  INV_X1    g0425(.A(new_n429), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n435), .A2(new_n437), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n625), .A2(new_n626), .B1(new_n442), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n305), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n309), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT89), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n560), .A2(new_n632), .ZN(new_n633));
  OAI221_X1 g0433(.A(KEYINPUT89), .B1(new_n265), .B2(new_n453), .C1(new_n260), .C2(new_n559), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n563), .A2(new_n260), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n306), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n572), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n640), .A3(G200), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n633), .A2(new_n634), .B1(new_n260), .B2(new_n563), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT90), .B1(new_n642), .B2(new_n335), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n567), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n461), .B1(new_n542), .B2(new_n497), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n527), .A2(new_n531), .A3(new_n534), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n545), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n639), .B1(new_n648), .B2(new_n621), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n639), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n614), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n567), .A2(new_n569), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n572), .A2(new_n573), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n615), .B2(new_n618), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n657), .B2(new_n652), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n448), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n631), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT91), .Z(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n488), .B2(new_n498), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n499), .A2(new_n669), .A3(new_n545), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n646), .A2(new_n668), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n668), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n529), .ZN(new_n676));
  MUX2_X1   g0476(.A(new_n538), .B(new_n647), .S(new_n676), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n647), .A2(new_n675), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n671), .A2(new_n681), .B1(new_n646), .B2(new_n675), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n211), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n548), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n218), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n644), .A2(new_n567), .B1(new_n572), .B2(new_n638), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n613), .A3(new_n596), .A4(new_n616), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT95), .B1(new_n692), .B2(new_n652), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n651), .A2(new_n694), .A3(KEYINPUT26), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(KEYINPUT29), .B(new_n675), .C1(new_n698), .C2(new_n649), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n675), .B1(new_n649), .B2(new_n658), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n457), .A2(new_n564), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n608), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n520), .A2(new_n525), .A3(new_n707), .A4(G179), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n709), .A3(KEYINPUT30), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT30), .B1(new_n705), .B2(new_n709), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n608), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n459), .A2(new_n637), .A3(new_n376), .A4(new_n526), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n713), .B2(new_n711), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n675), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n622), .A2(new_n675), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(KEYINPUT31), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n713), .A2(new_n718), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n723), .B(new_n675), .C1(new_n724), .C2(new_n710), .ZN(new_n725));
  OAI21_X1  g0525(.A(G330), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n703), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n690), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n291), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n207), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n685), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n214), .B1(G20), .B2(new_n306), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT98), .B(G159), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G20), .A3(new_n389), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT32), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n208), .A2(new_n376), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n389), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n201), .A2(new_n747), .B1(new_n749), .B2(new_n203), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(G179), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n208), .B1(new_n739), .B2(G190), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n546), .B1(new_n753), .B2(new_n501), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n389), .A3(G200), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n250), .B1(new_n755), .B2(new_n315), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n743), .A2(new_n750), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n744), .A2(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n744), .A2(KEYINPUT96), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(G190), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(new_n389), .A3(new_n760), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n757), .B1(new_n202), .B2(new_n761), .C1(new_n766), .C2(new_n343), .ZN(new_n767));
  XOR2_X1   g0567(.A(KEYINPUT33), .B(G317), .Z(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n749), .A2(new_n768), .B1(new_n755), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n747), .A2(new_n771), .B1(new_n753), .B2(new_n451), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n250), .B1(new_n741), .B2(G329), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n523), .B2(new_n752), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n770), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n761), .C1(new_n766), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n736), .B1(new_n767), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n735), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n211), .A2(G355), .A3(new_n250), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n684), .A2(new_n250), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n218), .ZN(new_n786));
  INV_X1    g0586(.A(G45), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n241), .A2(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n784), .B1(G116), .B2(new_n211), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n734), .B(new_n779), .C1(new_n783), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  INV_X1    g0591(.A(new_n782), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n677), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n679), .A2(new_n733), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G330), .B2(new_n677), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n735), .A2(new_n780), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n734), .B1(new_n343), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n334), .A2(new_n668), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n339), .B1(new_n331), .B2(new_n675), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n334), .ZN(new_n802));
  INV_X1    g0602(.A(new_n755), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n746), .A2(G303), .B1(new_n803), .B2(G87), .ZN(new_n804));
  INV_X1    g0604(.A(new_n753), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G97), .B1(new_n741), .B2(G311), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n256), .B1(new_n752), .B2(new_n315), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n806), .C1(KEYINPUT101), .C2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n748), .A2(KEYINPUT100), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G283), .B1(KEYINPUT101), .B2(new_n807), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n451), .B2(new_n761), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n808), .B(new_n814), .C1(G116), .C2(new_n765), .ZN(new_n815));
  INV_X1    g0615(.A(new_n761), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G143), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n747), .C1(new_n819), .C2(new_n749), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n765), .B2(new_n738), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n755), .A2(new_n203), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n250), .B1(new_n740), .B2(new_n825), .C1(new_n202), .C2(new_n753), .ZN(new_n826));
  INV_X1    g0626(.A(new_n752), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n824), .B(new_n826), .C1(G50), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n815), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n799), .B1(new_n781), .B2(new_n802), .C1(new_n829), .C2(new_n736), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n700), .B(new_n802), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n726), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n734), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n726), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(G384));
  NAND2_X1  g0636(.A1(new_n602), .A2(KEYINPUT35), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n216), .A2(new_n504), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(KEYINPUT35), .B2(new_n602), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n839), .B2(KEYINPUT103), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(KEYINPUT103), .B2(new_n839), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT36), .ZN(new_n842));
  INV_X1    g0642(.A(new_n218), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n207), .B(G13), .C1(new_n844), .C2(new_n237), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n666), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n430), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n435), .A2(new_n848), .A3(new_n425), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n435), .A2(new_n848), .A3(new_n851), .A4(new_n425), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(KEYINPUT38), .B(new_n853), .C1(new_n443), .C2(new_n848), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n848), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n438), .A2(new_n440), .B1(KEYINPUT18), .B2(new_n439), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n429), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n859), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n853), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n853), .B1(new_n443), .B2(new_n848), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n675), .B(new_n802), .C1(new_n649), .C2(new_n658), .ZN(new_n865));
  INV_X1    g0665(.A(new_n800), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n357), .A2(new_n675), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n386), .A2(new_n395), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n383), .B2(new_n385), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n864), .A2(new_n867), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n627), .A2(new_n442), .ZN(new_n875));
  INV_X1    g0675(.A(new_n853), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n848), .B1(new_n626), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n862), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n854), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(KEYINPUT39), .B2(new_n864), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n386), .A2(new_n675), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n874), .B1(new_n875), .B2(new_n847), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n448), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT105), .B1(new_n703), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n699), .A2(new_n448), .A3(new_n886), .A4(new_n702), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n631), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n883), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n802), .B1(new_n869), .B2(new_n871), .ZN(new_n891));
  INV_X1    g0691(.A(new_n720), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n575), .A2(new_n621), .A3(new_n668), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n723), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n705), .A2(new_n709), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT30), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n711), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n718), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n713), .B1(new_n711), .B2(new_n710), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT31), .B(new_n668), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT106), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT106), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n720), .A2(new_n903), .A3(KEYINPUT31), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n891), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n864), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n878), .B2(new_n854), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(new_n908), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n894), .A2(new_n905), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n448), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n448), .B2(new_n911), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n890), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n207), .B2(new_n730), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n890), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n846), .B1(new_n917), .B2(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n785), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n783), .B1(new_n211), .B2(new_n320), .C1(new_n920), .C2(new_n235), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n733), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n558), .A2(new_n566), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n668), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n639), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n691), .B2(new_n924), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(G317), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n256), .B1(new_n740), .B2(new_n928), .C1(new_n755), .C2(new_n501), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n747), .A2(new_n777), .B1(new_n753), .B2(new_n315), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(G303), .C2(new_n816), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT46), .B1(new_n752), .B2(new_n504), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n504), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n812), .A2(G294), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n931), .B(new_n934), .C1(new_n766), .C2(new_n769), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n746), .A2(G143), .B1(G137), .B2(new_n741), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n202), .B2(new_n752), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n812), .B2(new_n738), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n755), .A2(new_n343), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n256), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT111), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n938), .B(new_n941), .C1(new_n766), .C2(new_n201), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n753), .A2(new_n203), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n816), .B2(G150), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT110), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n935), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  OAI221_X1 g0747(.A(new_n922), .B1(new_n792), .B2(new_n927), .C1(new_n947), .C2(new_n736), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n671), .A2(new_n681), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n675), .A2(new_n606), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n621), .A2(new_n951), .B1(new_n614), .B2(new_n675), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT42), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n615), .A2(new_n618), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n952), .B(KEYINPUT107), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n957), .B2(new_n646), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n668), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n927), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n926), .B1(new_n960), .B2(KEYINPUT108), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT43), .B1(new_n962), .B2(new_n963), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n967), .A2(new_n968), .B1(new_n680), .B2(new_n956), .ZN(new_n969));
  INV_X1    g0769(.A(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n680), .A2(new_n956), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n971), .A3(new_n966), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n674), .A2(new_n681), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n950), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n679), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n727), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  INV_X1    g0778(.A(new_n680), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n682), .A2(new_n952), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT45), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n682), .A2(new_n952), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n978), .B(new_n979), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n978), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n981), .A2(new_n985), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n977), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n728), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n685), .B(KEYINPUT41), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n732), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n948), .B1(new_n973), .B2(new_n992), .ZN(G387));
  INV_X1    g0793(.A(new_n976), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n674), .A2(new_n792), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n232), .A2(new_n787), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT112), .Z(new_n997));
  OAI211_X1 g0797(.A(new_n687), .B(new_n787), .C1(new_n203), .C2(new_n343), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n323), .A2(new_n201), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n785), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n211), .A2(new_n250), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1004), .A2(new_n687), .B1(G107), .B2(new_n211), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n783), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n733), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n765), .A2(G68), .B1(new_n286), .B2(new_n748), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT114), .Z(new_n1009));
  OAI221_X1 g0809(.A(new_n250), .B1(new_n740), .B2(new_n819), .C1(new_n755), .C2(new_n501), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n746), .A2(G159), .B1(new_n570), .B2(new_n805), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n343), .B2(new_n752), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G50), .C2(new_n816), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n752), .A2(new_n451), .B1(new_n753), .B2(new_n769), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n816), .A2(G317), .B1(G322), .B2(new_n746), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n777), .B2(new_n811), .C1(new_n766), .C2(new_n523), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT115), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1018), .B2(KEYINPUT48), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT48), .B2(new_n1018), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n256), .B1(new_n740), .B2(new_n771), .C1(new_n755), .C2(new_n504), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT116), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1014), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1007), .B1(new_n1026), .B2(new_n735), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n994), .A2(new_n732), .B1(new_n995), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n977), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(KEYINPUT117), .A3(new_n685), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n728), .B2(new_n994), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT117), .B1(new_n1029), .B2(new_n685), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  OR3_X1    g0833(.A1(new_n984), .A2(new_n988), .A3(new_n977), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n685), .A3(new_n989), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n732), .B1(new_n984), .B2(new_n988), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n256), .B1(new_n741), .B2(G143), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n203), .B2(new_n752), .C1(new_n469), .C2(new_n755), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT118), .Z(new_n1039));
  INV_X1    g0839(.A(G159), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n1040), .B1(new_n819), .B2(new_n747), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT51), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n765), .A2(new_n323), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n753), .A2(new_n343), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n812), .B2(G50), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT119), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n761), .A2(new_n777), .B1(new_n928), .B2(new_n747), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT52), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n256), .B1(new_n740), .B2(new_n776), .C1(new_n755), .C2(new_n315), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n752), .A2(new_n769), .B1(new_n753), .B2(new_n504), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n812), .C2(G303), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n451), .B2(new_n766), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1048), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n735), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n785), .A2(new_n244), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n735), .B(new_n782), .C1(new_n684), .C2(G97), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n734), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(new_n957), .C2(new_n792), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1035), .A2(new_n1036), .A3(new_n1061), .ZN(G390));
  NAND2_X1  g0862(.A1(new_n906), .A2(G330), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT39), .ZN(new_n1065));
  AOI21_X1  g0865(.A(KEYINPUT38), .B1(new_n859), .B2(new_n853), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n855), .B2(new_n854), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1065), .B1(new_n1067), .B2(new_n860), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n882), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n867), .B2(new_n873), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1068), .A2(new_n1070), .A3(new_n880), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n879), .A2(new_n882), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n649), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n693), .B(new_n695), .C1(KEYINPUT26), .C2(new_n657), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n668), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n801), .A2(new_n334), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n800), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1072), .B1(new_n1078), .B2(new_n873), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1064), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n802), .C1(new_n722), .C2(new_n725), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(new_n872), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n882), .B(new_n879), .C1(new_n1077), .C2(new_n872), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n881), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1083), .C1(new_n1084), .C2(new_n1070), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G330), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n894), .B2(new_n905), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1088), .A2(new_n448), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n630), .B(new_n1089), .C1(new_n885), .C2(new_n887), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1081), .A2(new_n872), .B1(G330), .B2(new_n906), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n867), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1077), .B1(new_n1081), .B2(new_n872), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n873), .B1(new_n1088), .B2(new_n802), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1086), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1080), .A2(new_n1090), .A3(new_n1085), .A4(new_n1095), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n685), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1080), .A2(new_n732), .A3(new_n1085), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n798), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n733), .B1(new_n286), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n812), .A2(G137), .B1(G132), .B2(new_n816), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n250), .B1(new_n740), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n755), .A2(new_n201), .B1(new_n753), .B2(new_n1040), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G128), .C2(new_n746), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n752), .A2(new_n819), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1103), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n766), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n812), .A2(G107), .B1(G116), .B2(new_n816), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n250), .B(new_n824), .C1(G294), .C2(new_n741), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n752), .A2(new_n469), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1044), .B(new_n1115), .C1(G283), .C2(new_n746), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n766), .A2(new_n501), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1110), .A2(new_n1112), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1102), .B1(new_n1119), .B2(new_n735), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1084), .B2(new_n781), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1100), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1099), .A2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n907), .A2(new_n908), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n906), .A2(new_n909), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(G330), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT122), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(KEYINPUT122), .A3(G330), .A4(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n305), .A2(new_n309), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n308), .A2(new_n847), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1135), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1129), .A2(new_n1130), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n883), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1127), .A2(new_n1128), .A3(new_n1139), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1124), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1098), .A2(new_n1090), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1130), .A2(new_n1140), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT122), .B1(new_n910), .B2(G330), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1143), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n883), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(KEYINPUT123), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1146), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1152), .A2(new_n1147), .A3(KEYINPUT57), .A4(new_n1153), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n685), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1146), .A2(new_n732), .A3(new_n1154), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n749), .A2(new_n825), .B1(new_n752), .B2(new_n1111), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n746), .A2(G125), .B1(G150), .B2(new_n805), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G128), .C2(new_n816), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n766), .B2(new_n818), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n803), .A2(new_n738), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n741), .C2(G124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n501), .A2(new_n749), .B1(new_n747), .B2(new_n504), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n202), .A2(new_n755), .B1(new_n752), .B2(new_n343), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n256), .B(new_n267), .C1(new_n740), .C2(new_n769), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n943), .A4(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n315), .B2(new_n761), .C1(new_n766), .C2(new_n320), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n201), .B1(new_n254), .B2(G41), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n1172), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n733), .B1(G50), .B2(new_n1101), .C1(new_n1182), .C2(new_n736), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1140), .B2(new_n780), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT121), .Z(new_n1185));
  NAND2_X1  g0985(.A1(new_n1162), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1161), .A2(new_n1187), .ZN(G375));
  NOR2_X1   g0988(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1081), .A2(new_n872), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1092), .B1(new_n1190), .B2(new_n1063), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1089), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n888), .A2(new_n631), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1096), .A3(new_n991), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n811), .A2(new_n504), .B1(new_n769), .B2(new_n761), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n250), .B(new_n939), .C1(G303), .C2(new_n741), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n827), .A2(G97), .B1(new_n805), .B2(new_n570), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n451), .C2(new_n747), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(G107), .C2(new_n765), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n811), .A2(new_n1111), .B1(new_n818), .B2(new_n761), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n755), .A2(new_n202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n256), .B(new_n1203), .C1(G128), .C2(new_n741), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n746), .A2(G132), .B1(G50), .B2(new_n805), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1040), .C2(new_n752), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1202), .B(new_n1206), .C1(G150), .C2(new_n765), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n735), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n733), .C1(G68), .C2(new_n1101), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n872), .B2(new_n780), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1095), .B2(new_n732), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1196), .A2(new_n1211), .ZN(G381));
  INV_X1    g1012(.A(G390), .ZN(new_n1213));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G396), .A2(new_n1215), .A3(G393), .A4(G381), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1216), .A2(G387), .A3(new_n1218), .ZN(G407));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  OAI21_X1  g1020(.A(KEYINPUT60), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(new_n1195), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1192), .A2(KEYINPUT60), .A3(new_n1194), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n685), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1211), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1214), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G384), .B(new_n1211), .C1(new_n1222), .C2(new_n1224), .ZN(new_n1227));
  INV_X1    g1027(.A(G2897), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n667), .A2(G213), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1226), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1228), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1221), .A2(new_n1195), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n685), .A3(new_n1223), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G384), .B1(new_n1234), .B2(new_n1211), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1231), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1159), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1238));
  OAI21_X1  g1038(.A(G378), .B1(new_n1238), .B2(new_n1186), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1152), .A2(new_n732), .A3(new_n1153), .ZN(new_n1240));
  AND4_X1   g1040(.A1(new_n1099), .A2(new_n1240), .A3(new_n1122), .A4(new_n1185), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1146), .A2(new_n991), .A3(new_n1154), .A4(new_n1147), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1241), .A2(new_n1242), .B1(G213), .B2(new_n667), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1237), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT126), .B1(new_n1244), .B2(KEYINPUT61), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1239), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT62), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1239), .A2(KEYINPUT124), .A3(new_n1243), .A4(new_n1246), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1229), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G375), .B2(G378), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1256), .B(new_n1257), .C1(new_n1260), .C2(new_n1237), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1249), .A2(KEYINPUT127), .A3(new_n1255), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1213), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(G396), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G390), .B(new_n948), .C1(new_n973), .C2(new_n992), .ZN(new_n1270));
  AND4_X1   g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(KEYINPUT125), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1272), .A2(new_n1269), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(new_n1266), .A3(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1274), .A2(KEYINPUT61), .A3(new_n1244), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1246), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(KEYINPUT63), .C2(new_n1253), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(G405));
  NAND2_X1  g1079(.A1(new_n1218), .A2(new_n1239), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1246), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1274), .ZN(G402));
endmodule


