//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OR3_X1    g004(.A1(new_n204), .A2(KEYINPUT26), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT27), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT27), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT66), .B1(new_n213), .B2(G183gat), .ZN(new_n217));
  AOI21_X1  g016(.A(G190gat), .B1(new_n213), .B2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(new_n211), .A3(KEYINPUT27), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n215), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n216), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT23), .B1(new_n205), .B2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n228), .B(new_n229), .C1(G169gat), .C2(G176gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(new_n202), .C2(new_n203), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n210), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n233), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n204), .B1(KEYINPUT23), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n207), .A2(new_n235), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n238), .A3(new_n239), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(new_n230), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n232), .A2(new_n241), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n226), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n254), .B2(new_n253), .ZN(new_n256));
  XOR2_X1   g055(.A(G127gat), .B(G134gat), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n250), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n248), .B(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT32), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  XOR2_X1   g070(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G15gat), .B(G43gat), .Z(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n278), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(new_n272), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n271), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n279), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n269), .B(new_n270), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(KEYINPUT22), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n226), .B2(new_n247), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n234), .A2(new_n235), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n207), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n240), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n230), .A4(new_n243), .ZN(new_n303));
  INV_X1    g102(.A(new_n245), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n233), .B1(new_n231), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n221), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT67), .B1(new_n221), .B2(new_n215), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(new_n308), .A3(new_n216), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(KEYINPUT72), .C1(new_n309), .C2(new_n209), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n299), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(new_n312), .C1(new_n226), .C2(new_n247), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n297), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n310), .A3(new_n315), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n312), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n312), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT74), .B1(new_n248), .B2(new_n312), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n324), .B(new_n313), .C1(new_n226), .C2(new_n247), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n317), .B1(new_n327), .B2(new_n297), .ZN(new_n328));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  OAI21_X1  g130(.A(new_n289), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n319), .A2(new_n320), .B1(new_n323), .B2(new_n325), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n296), .B1(new_n334), .B2(new_n322), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT75), .B(new_n333), .C1(new_n335), .C2(new_n317), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n338));
  NOR4_X1   g137(.A1(new_n335), .A2(new_n338), .A3(new_n317), .A4(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT30), .B1(new_n328), .B2(new_n331), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n288), .A2(new_n337), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n339), .A2(new_n341), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n288), .B1(new_n344), .B2(new_n337), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n287), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G1gat), .B(G29gat), .Z(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  INV_X1    g154(.A(G155gat), .ZN(new_n356));
  INV_X1    g155(.A(G162gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(KEYINPUT2), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT78), .B(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G141gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n361), .A2(G148gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n358), .A2(KEYINPUT77), .A3(new_n355), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT77), .B1(new_n358), .B2(new_n355), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n258), .A3(new_n263), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n258), .B2(new_n263), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n354), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n373), .A2(new_n380), .A3(new_n258), .A4(new_n263), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n387), .A2(new_n264), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n354), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n378), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n379), .A2(new_n392), .A3(new_n381), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n374), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n391), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n352), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n389), .A2(new_n382), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n351), .B(new_n396), .C1(new_n399), .C2(new_n378), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT6), .B(new_n352), .C1(new_n390), .C2(new_n397), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n296), .A2(new_n315), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n373), .B1(new_n405), .B2(new_n386), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n315), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n297), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  INV_X1    g210(.A(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n410), .B(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n404), .A2(KEYINPUT35), .A3(new_n420), .ZN(new_n421));
  AOI211_X1 g220(.A(new_n333), .B(new_n317), .C1(new_n327), .C2(new_n297), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n332), .A2(new_n336), .B1(KEYINPUT30), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n271), .B1(new_n279), .B2(new_n281), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n283), .A2(new_n284), .ZN(new_n427));
  INV_X1    g226(.A(new_n420), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n341), .B1(new_n403), .B2(new_n402), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n425), .A2(new_n429), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n346), .A2(new_n421), .B1(new_n432), .B2(KEYINPUT35), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n423), .B2(new_n424), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n337), .A2(new_n424), .A3(new_n340), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n420), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT36), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n282), .B2(new_n285), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT36), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n354), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n443), .A2(new_n354), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  INV_X1    g246(.A(new_n376), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n374), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n354), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(KEYINPUT85), .A3(new_n374), .A4(new_n353), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT39), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n351), .B(new_n445), .C1(new_n446), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT86), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n446), .A2(new_n452), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n445), .A2(new_n351), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT40), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n398), .A2(KEYINPUT40), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n453), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n343), .B2(new_n345), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n331), .B1(new_n328), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n327), .A2(new_n296), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n314), .A2(new_n316), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n468), .B2(new_n297), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT38), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT87), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n328), .A2(new_n331), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n402), .A2(new_n474), .A3(new_n403), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n466), .B1(new_n465), .B2(new_n328), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(KEYINPUT38), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n420), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n441), .B1(new_n442), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n478), .A3(KEYINPUT88), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n433), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(G1gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT16), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n485), .B2(G1gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(KEYINPUT92), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT92), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n488), .B2(new_n491), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G43gat), .A2(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT90), .B(G50gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(G43gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(G43gat), .A2(G50gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT15), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n507), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n506), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n506), .A2(new_n511), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n512), .A2(new_n513), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT17), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n494), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n488), .A2(new_n491), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(KEYINPUT94), .A3(new_n515), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT95), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT18), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(KEYINPUT95), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n515), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT13), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n531), .A2(new_n537), .A3(new_n539), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n530), .A2(KEYINPUT18), .B1(new_n544), .B2(new_n543), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(KEYINPUT97), .A3(new_n537), .A4(new_n539), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n539), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n536), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT98), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n522), .B1(KEYINPUT21), .B2(new_n560), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n568), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT103), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n517), .B(new_n518), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n578), .B(new_n579), .Z(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT101), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n580), .A2(new_n588), .A3(new_n581), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT102), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT102), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n580), .A2(new_n585), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n594), .A2(new_n581), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n577), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n515), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n576), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n575), .A2(KEYINPUT103), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT99), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n603), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n576), .B(new_n609), .C1(new_n597), .C2(new_n601), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n604), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n604), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n595), .A2(new_n590), .A3(new_n560), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n618), .B(new_n619), .C1(new_n598), .C2(new_n560), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n560), .A2(KEYINPUT10), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n596), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n619), .ZN(new_n628));
  INV_X1    g427(.A(new_n560), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n596), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n625), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n617), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n626), .B(new_n616), .C1(new_n625), .C2(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n573), .A2(new_n613), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n482), .A2(new_n555), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n404), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g438(.A1(new_n343), .A2(new_n345), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n490), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(KEYINPUT42), .B2(new_n644), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n637), .A2(new_n648), .A3(new_n286), .ZN(new_n649));
  INV_X1    g448(.A(new_n440), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n637), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n651), .B2(new_n648), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n420), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n460), .A2(new_n462), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n344), .A2(new_n337), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT84), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n344), .A2(new_n288), .A3(new_n337), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n472), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n333), .B1(new_n335), .B2(new_n317), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n333), .A2(KEYINPUT37), .ZN(new_n665));
  INV_X1    g464(.A(new_n328), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(KEYINPUT37), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n404), .B(new_n474), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n428), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n442), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n441), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n481), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n346), .A2(new_n421), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n432), .A2(KEYINPUT35), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n613), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n573), .A2(new_n555), .A3(new_n634), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n504), .A3(new_n404), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n482), .B2(new_n613), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n676), .ZN(new_n684));
  INV_X1    g483(.A(new_n613), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n678), .ZN(new_n688));
  INV_X1    g487(.A(new_n404), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n681), .A2(new_n690), .ZN(G1328gat));
  OAI21_X1  g490(.A(G36gat), .B1(new_n688), .B2(new_n640), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n679), .A2(new_n505), .A3(new_n641), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n697), .B2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n650), .A3(new_n686), .A4(new_n678), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(G43gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n287), .A2(G43gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n677), .A2(new_n678), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n701), .B2(G43gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n700), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n701), .A2(G43gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n704), .A4(new_n703), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n687), .A2(new_n420), .A3(new_n678), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n498), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT107), .ZN(new_n720));
  INV_X1    g519(.A(new_n498), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n679), .A2(new_n420), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n719), .B(new_n722), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n573), .A2(new_n613), .A3(new_n634), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n482), .A2(new_n554), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n404), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n641), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n650), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n287), .A2(G71gat), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n736), .A2(G71gat), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n420), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n573), .A2(new_n554), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n635), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n687), .A2(new_n404), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n583), .B1(new_n745), .B2(KEYINPUT108), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT108), .B2(new_n745), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n677), .A2(KEYINPUT51), .A3(new_n742), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n677), .B2(new_n742), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n404), .A2(new_n583), .A3(new_n634), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT109), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n747), .B1(new_n750), .B2(new_n752), .ZN(G1336gat));
  NOR3_X1   g552(.A1(new_n640), .A2(G92gat), .A3(new_n635), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT111), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n748), .B2(new_n749), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT112), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n758), .B(new_n755), .C1(new_n748), .C2(new_n749), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n683), .A2(new_n641), .A3(new_n686), .A4(new_n744), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n757), .B(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  NAND2_X1  g563(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n762), .B(new_n765), .C1(new_n756), .C2(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  OR4_X1    g566(.A1(G99gat), .A2(new_n750), .A3(new_n287), .A4(new_n635), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n687), .A2(new_n650), .A3(new_n744), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G99gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n683), .A2(new_n420), .A3(new_n686), .A4(new_n744), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT113), .B1(new_n772), .B2(G106gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n428), .A2(G106gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n634), .B(new_n774), .C1(new_n748), .C2(new_n749), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n622), .B1(new_n630), .B2(new_n618), .ZN(new_n779));
  INV_X1    g578(.A(new_n625), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT54), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n624), .A2(new_n625), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n626), .A2(new_n784), .A3(KEYINPUT114), .A4(KEYINPUT54), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n617), .B1(new_n626), .B2(KEYINPUT54), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n633), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n787), .B1(new_n783), .B2(new_n785), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(KEYINPUT55), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n794), .A3(new_n554), .ZN(new_n795));
  INV_X1    g594(.A(new_n544), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n527), .A2(new_n541), .A3(new_n796), .A4(new_n542), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n577), .A2(new_n494), .B1(new_n525), .B2(new_n526), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n528), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n535), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT115), .Z(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n551), .A3(new_n634), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n685), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n613), .B1(new_n790), .B2(new_n789), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n801), .A2(new_n551), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(new_n794), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT116), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n805), .A3(new_n794), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n801), .A2(new_n551), .A3(new_n634), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n789), .A2(new_n790), .B1(new_n551), .B2(new_n553), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n794), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n685), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n807), .A2(new_n813), .A3(new_n572), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n636), .A2(new_n554), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n420), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n817), .A2(new_n404), .A3(new_n346), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n554), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n634), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n573), .ZN(new_n823));
  NOR2_X1   g622(.A1(KEYINPUT117), .A2(G127gat), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n823), .B(new_n824), .Z(G1342gat));
  AOI21_X1  g624(.A(new_n613), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n827), .B(new_n828), .Z(G1343gat));
  NAND2_X1  g628(.A1(new_n795), .A2(new_n802), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n613), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT119), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n803), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n809), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n815), .B1(new_n835), .B2(new_n572), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT57), .B1(new_n836), .B2(new_n428), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n814), .A2(new_n816), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n420), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n641), .A2(new_n650), .A3(new_n689), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT118), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n555), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n838), .A2(new_n420), .A3(new_n841), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n555), .A2(G141gat), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT58), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n840), .A2(new_n842), .ZN(new_n849));
  INV_X1    g648(.A(new_n834), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n809), .B1(new_n803), .B2(new_n833), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n572), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n816), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n839), .B1(new_n853), .B2(new_n420), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n856), .A3(new_n840), .A4(new_n842), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n554), .A3(new_n857), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n858), .A2(G141gat), .B1(new_n845), .B2(new_n846), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n848), .B1(new_n859), .B2(new_n860), .ZN(G1344gat));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n855), .A2(new_n634), .A3(new_n857), .ZN(new_n863));
  INV_X1    g662(.A(new_n360), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n839), .B(new_n428), .C1(new_n814), .C2(new_n816), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n573), .B1(new_n831), .B2(new_n809), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n420), .B1(new_n869), .B2(new_n815), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT121), .B1(new_n870), .B2(new_n839), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n634), .A3(new_n842), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n862), .A2(new_n363), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n635), .A2(new_n360), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n873), .A2(new_n874), .B1(new_n845), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n865), .A2(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n845), .A2(new_n356), .A3(new_n573), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n855), .A2(new_n573), .A3(new_n857), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n356), .ZN(G1346gat));
  NAND3_X1  g679(.A1(new_n855), .A2(new_n685), .A3(new_n857), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT122), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n855), .A2(new_n883), .A3(new_n685), .A4(new_n857), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(G162gat), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n845), .A2(new_n357), .A3(new_n685), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n640), .A2(new_n404), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n838), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(new_n429), .ZN(new_n890));
  AOI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n554), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n888), .B(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n286), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT124), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(KEYINPUT124), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n817), .A3(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n202), .A3(new_n555), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n891), .A2(new_n897), .ZN(G1348gat));
  OAI21_X1  g697(.A(G176gat), .B1(new_n896), .B2(new_n635), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n890), .A2(new_n203), .A3(new_n634), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  NOR2_X1   g700(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n572), .A2(new_n214), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT125), .B1(new_n890), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n896), .B2(new_n572), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n210), .A3(new_n685), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n896), .A2(new_n613), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n911), .A2(new_n210), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n911), .B2(new_n210), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(G1351gat));
  AND3_X1   g714(.A1(new_n889), .A2(new_n420), .A3(new_n440), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n554), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n892), .A2(new_n440), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n872), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n554), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(new_n634), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n925));
  OAI21_X1  g724(.A(G204gat), .B1(new_n919), .B2(new_n635), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n916), .A2(new_n291), .A3(new_n573), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n872), .A2(new_n573), .A3(new_n918), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n919), .B2(new_n613), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n292), .A3(new_n685), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


