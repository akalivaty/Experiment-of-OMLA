

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758;

  XNOR2_X1 U368 ( .A(n393), .B(n361), .ZN(n758) );
  XNOR2_X1 U369 ( .A(n417), .B(n360), .ZN(n422) );
  NOR2_X1 U370 ( .A1(n674), .A2(n673), .ZN(n410) );
  XNOR2_X1 U371 ( .A(n349), .B(n444), .ZN(n369) );
  NOR2_X2 U372 ( .A1(n428), .A2(n425), .ZN(n368) );
  NOR2_X2 U373 ( .A1(n601), .A2(n355), .ZN(n603) );
  OR2_X2 U374 ( .A1(n717), .A2(G902), .ZN(n395) );
  NAND2_X1 U375 ( .A1(n346), .A2(n359), .ZN(n399) );
  NAND2_X1 U376 ( .A1(n402), .A2(n401), .ZN(n346) );
  NOR2_X1 U377 ( .A1(n681), .A2(n680), .ZN(n684) );
  NAND2_X1 U378 ( .A1(n579), .A2(n684), .ZN(n607) );
  AND2_X2 U379 ( .A1(n666), .A2(n628), .ZN(n629) );
  NOR2_X2 U380 ( .A1(n437), .A2(n560), .ZN(n364) );
  NAND2_X1 U381 ( .A1(n629), .A2(n665), .ZN(n413) );
  AND2_X1 U382 ( .A1(n378), .A2(n387), .ZN(n384) );
  NOR2_X1 U383 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U384 ( .A1(n614), .A2(n650), .ZN(n616) );
  AND2_X1 U385 ( .A1(n377), .A2(n376), .ZN(n385) );
  NAND2_X1 U386 ( .A1(n415), .A2(n397), .ZN(n389) );
  AND2_X1 U387 ( .A1(n577), .A2(n579), .ZN(n590) );
  XNOR2_X1 U388 ( .A(n596), .B(KEYINPUT38), .ZN(n671) );
  INV_X1 U389 ( .A(n578), .ZN(n596) );
  XNOR2_X1 U390 ( .A(n608), .B(KEYINPUT6), .ZN(n565) );
  OR2_X1 U391 ( .A1(n568), .A2(n587), .ZN(n673) );
  XNOR2_X1 U392 ( .A(n395), .B(n465), .ZN(n576) );
  INV_X2 U393 ( .A(G953), .ZN(n735) );
  NOR2_X1 U394 ( .A1(n714), .A2(n729), .ZN(n715) );
  XNOR2_X1 U395 ( .A(n720), .B(n347), .ZN(n721) );
  XOR2_X1 U396 ( .A(n719), .B(n718), .Z(n347) );
  BUF_X1 U397 ( .A(n716), .Z(n725) );
  XNOR2_X1 U398 ( .A(n713), .B(n712), .ZN(n714) );
  BUF_X1 U399 ( .A(n666), .Z(n348) );
  XNOR2_X1 U400 ( .A(n743), .B(G101), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n743), .B(G101), .ZN(n438) );
  XNOR2_X1 U402 ( .A(n438), .B(n542), .ZN(n414) );
  XNOR2_X1 U403 ( .A(n742), .B(G146), .ZN(n444) );
  XNOR2_X1 U404 ( .A(n437), .B(n409), .ZN(n567) );
  INV_X1 U405 ( .A(KEYINPUT94), .ZN(n409) );
  INV_X1 U406 ( .A(KEYINPUT83), .ZN(n375) );
  OR2_X1 U407 ( .A1(n660), .A2(n675), .ZN(n376) );
  XNOR2_X1 U408 ( .A(G116), .B(G113), .ZN(n498) );
  INV_X1 U409 ( .A(G128), .ZN(n458) );
  XNOR2_X1 U410 ( .A(n540), .B(n468), .ZN(n514) );
  XNOR2_X1 U411 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n468) );
  XOR2_X1 U412 ( .A(G137), .B(G140), .Z(n515) );
  XNOR2_X1 U413 ( .A(KEYINPUT92), .B(G110), .ZN(n460) );
  XNOR2_X1 U414 ( .A(n419), .B(n457), .ZN(n580) );
  INV_X1 U415 ( .A(G478), .ZN(n440) );
  XNOR2_X1 U416 ( .A(n522), .B(n521), .ZN(n681) );
  XNOR2_X1 U417 ( .A(G119), .B(G128), .ZN(n508) );
  XOR2_X1 U418 ( .A(G122), .B(G107), .Z(n486) );
  XNOR2_X1 U419 ( .A(n492), .B(n352), .ZN(n443) );
  XOR2_X1 U420 ( .A(KEYINPUT99), .B(G140), .Z(n474) );
  XNOR2_X1 U421 ( .A(n410), .B(n418), .ZN(n701) );
  INV_X1 U422 ( .A(KEYINPUT41), .ZN(n418) );
  XNOR2_X1 U423 ( .A(n555), .B(KEYINPUT67), .ZN(n556) );
  BUF_X1 U424 ( .A(n466), .Z(n683) );
  AND2_X1 U425 ( .A1(n589), .A2(n375), .ZN(n373) );
  INV_X1 U426 ( .A(n575), .ZN(n396) );
  XNOR2_X1 U427 ( .A(KEYINPUT76), .B(KEYINPUT5), .ZN(n501) );
  XOR2_X1 U428 ( .A(G137), .B(KEYINPUT98), .Z(n502) );
  XNOR2_X1 U429 ( .A(n469), .B(n445), .ZN(n742) );
  INV_X1 U430 ( .A(G134), .ZN(n445) );
  XNOR2_X1 U431 ( .A(n446), .B(KEYINPUT70), .ZN(n469) );
  INV_X1 U432 ( .A(G131), .ZN(n446) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n475) );
  XOR2_X1 U434 ( .A(G143), .B(G122), .Z(n473) );
  XNOR2_X1 U435 ( .A(n500), .B(n499), .ZN(n547) );
  XOR2_X1 U436 ( .A(KEYINPUT3), .B(G119), .Z(n499) );
  INV_X1 U437 ( .A(KEYINPUT71), .ZN(n497) );
  NAND2_X1 U438 ( .A1(n453), .A2(KEYINPUT82), .ZN(n452) );
  XNOR2_X1 U439 ( .A(KEYINPUT15), .B(G902), .ZN(n627) );
  INV_X1 U440 ( .A(G237), .ZN(n533) );
  XNOR2_X1 U441 ( .A(n566), .B(KEYINPUT33), .ZN(n669) );
  NAND2_X1 U442 ( .A1(n609), .A2(n573), .ZN(n566) );
  INV_X1 U443 ( .A(G902), .ZN(n534) );
  XNOR2_X1 U444 ( .A(n576), .B(n448), .ZN(n466) );
  INV_X1 U445 ( .A(KEYINPUT1), .ZN(n448) );
  XNOR2_X1 U446 ( .A(n369), .B(n464), .ZN(n717) );
  INV_X1 U447 ( .A(G146), .ZN(n467) );
  XNOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n538) );
  NAND2_X1 U449 ( .A1(n701), .A2(n590), .ZN(n417) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT39), .ZN(n604) );
  INV_X1 U451 ( .A(n583), .ZN(n391) );
  NOR2_X1 U452 ( .A1(n596), .A2(n350), .ZN(n433) );
  INV_X1 U453 ( .A(n608), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n405), .B(KEYINPUT97), .ZN(n439) );
  INV_X1 U455 ( .A(n607), .ZN(n408) );
  XNOR2_X1 U456 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U457 ( .A(n442), .B(n441), .ZN(n722) );
  XNOR2_X1 U458 ( .A(n493), .B(n495), .ZN(n441) );
  XNOR2_X1 U459 ( .A(n443), .B(n494), .ZN(n442) );
  XNOR2_X1 U460 ( .A(n482), .B(n481), .ZN(n632) );
  XNOR2_X1 U461 ( .A(n480), .B(n456), .ZN(n481) );
  AND2_X1 U462 ( .A1(n635), .A2(G953), .ZN(n729) );
  INV_X1 U463 ( .A(KEYINPUT32), .ZN(n454) );
  XNOR2_X1 U464 ( .A(n610), .B(KEYINPUT31), .ZN(n660) );
  AND2_X1 U465 ( .A1(n611), .A2(n447), .ZN(n612) );
  NAND2_X1 U466 ( .A1(n439), .A2(n398), .ZN(n647) );
  XOR2_X1 U467 ( .A(KEYINPUT81), .B(n529), .Z(n350) );
  AND2_X1 U468 ( .A1(n608), .A2(n396), .ZN(n351) );
  XNOR2_X1 U469 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n352) );
  AND2_X1 U470 ( .A1(n391), .A2(n390), .ZN(n353) );
  AND2_X1 U471 ( .A1(n587), .A2(n568), .ZN(n354) );
  NOR2_X1 U472 ( .A1(n600), .A2(n447), .ZN(n355) );
  AND2_X1 U473 ( .A1(n548), .A2(G210), .ZN(n356) );
  INV_X1 U474 ( .A(n675), .ZN(n411) );
  NAND2_X1 U475 ( .A1(n594), .A2(n595), .ZN(n357) );
  AND2_X1 U476 ( .A1(n411), .A2(n398), .ZN(n358) );
  NAND2_X1 U477 ( .A1(n616), .A2(KEYINPUT44), .ZN(n359) );
  XNOR2_X1 U478 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n360) );
  XOR2_X1 U479 ( .A(n584), .B(KEYINPUT40), .Z(n361) );
  XOR2_X1 U480 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n362) );
  XNOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n363) );
  INV_X1 U482 ( .A(KEYINPUT88), .ZN(n406) );
  XNOR2_X1 U483 ( .A(n414), .B(n736), .ZN(n709) );
  BUF_X1 U484 ( .A(n615), .Z(n367) );
  XNOR2_X1 U485 ( .A(n455), .B(n454), .ZN(n614) );
  NAND2_X1 U486 ( .A1(n385), .A2(n389), .ZN(n379) );
  XNOR2_X1 U487 ( .A(n364), .B(KEYINPUT22), .ZN(n613) );
  XNOR2_X2 U488 ( .A(n365), .B(KEYINPUT110), .ZN(n757) );
  NAND2_X1 U489 ( .A1(n434), .A2(n354), .ZN(n365) );
  XNOR2_X2 U490 ( .A(n366), .B(n363), .ZN(n730) );
  NAND2_X1 U491 ( .A1(n404), .A2(n399), .ZN(n366) );
  NAND2_X1 U492 ( .A1(n368), .A2(n431), .ZN(n601) );
  XNOR2_X1 U493 ( .A(n369), .B(n420), .ZN(n638) );
  INV_X1 U494 ( .A(n432), .ZN(n374) );
  NAND2_X1 U495 ( .A1(n371), .A2(n370), .ZN(n432) );
  NAND2_X1 U496 ( .A1(n373), .A2(n757), .ZN(n370) );
  NAND2_X1 U497 ( .A1(n372), .A2(KEYINPUT83), .ZN(n371) );
  NAND2_X1 U498 ( .A1(n757), .A2(n589), .ZN(n372) );
  NAND2_X1 U499 ( .A1(n374), .A2(n595), .ZN(n424) );
  NAND2_X1 U500 ( .A1(n439), .A2(n358), .ZN(n377) );
  NAND2_X1 U501 ( .A1(n379), .A2(n406), .ZN(n378) );
  NAND2_X1 U502 ( .A1(n380), .A2(n388), .ZN(n383) );
  NAND2_X1 U503 ( .A1(n389), .A2(KEYINPUT88), .ZN(n381) );
  INV_X1 U504 ( .A(n385), .ZN(n382) );
  NAND2_X1 U505 ( .A1(n384), .A2(n383), .ZN(n404) );
  NAND2_X1 U506 ( .A1(n615), .A2(KEYINPUT44), .ZN(n388) );
  NAND2_X1 U507 ( .A1(n615), .A2(n386), .ZN(n387) );
  AND2_X1 U508 ( .A1(n406), .A2(KEYINPUT44), .ZN(n386) );
  XNOR2_X2 U509 ( .A(n571), .B(n570), .ZN(n615) );
  XNOR2_X2 U510 ( .A(n564), .B(KEYINPUT75), .ZN(n609) );
  NAND2_X1 U511 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U512 ( .A1(n669), .A2(n567), .ZN(n412) );
  NAND2_X1 U513 ( .A1(n616), .A2(n403), .ZN(n402) );
  NAND2_X1 U514 ( .A1(n407), .A2(n554), .ZN(n557) );
  XNOR2_X1 U515 ( .A(n389), .B(G101), .ZN(G3) );
  NOR2_X1 U516 ( .A1(n607), .A2(n350), .ZN(n390) );
  NOR2_X1 U517 ( .A1(n583), .A2(n607), .ZN(n392) );
  AND2_X1 U518 ( .A1(n392), .A2(n433), .ZN(n436) );
  NAND2_X1 U519 ( .A1(n604), .A2(n655), .ZN(n393) );
  NAND2_X1 U520 ( .A1(n353), .A2(n671), .ZN(n394) );
  NAND2_X1 U521 ( .A1(n466), .A2(n684), .ZN(n564) );
  NOR2_X1 U522 ( .A1(n608), .A2(n397), .ZN(n611) );
  INV_X1 U523 ( .A(n681), .ZN(n397) );
  NAND2_X1 U524 ( .A1(n688), .A2(n398), .ZN(n689) );
  INV_X1 U525 ( .A(KEYINPUT44), .ZN(n401) );
  INV_X1 U526 ( .A(n615), .ZN(n403) );
  NAND2_X1 U527 ( .A1(n567), .A2(n408), .ZN(n405) );
  XNOR2_X2 U528 ( .A(n557), .B(n556), .ZN(n437) );
  NAND2_X1 U529 ( .A1(n590), .A2(n407), .ZN(n591) );
  XNOR2_X2 U530 ( .A(n551), .B(KEYINPUT19), .ZN(n407) );
  XNOR2_X1 U531 ( .A(n416), .B(KEYINPUT87), .ZN(n415) );
  XNOR2_X1 U532 ( .A(n412), .B(n362), .ZN(n449) );
  XNOR2_X2 U533 ( .A(n413), .B(n630), .ZN(n716) );
  BUF_X2 U534 ( .A(n580), .Z(n608) );
  NAND2_X1 U535 ( .A1(n709), .A2(n627), .ZN(n549) );
  NAND2_X1 U536 ( .A1(n613), .A2(n574), .ZN(n416) );
  INV_X1 U537 ( .A(n422), .ZN(n756) );
  NAND2_X1 U538 ( .A1(n638), .A2(n534), .ZN(n419) );
  XNOR2_X1 U539 ( .A(n506), .B(n505), .ZN(n420) );
  NAND2_X1 U540 ( .A1(n422), .A2(n421), .ZN(n430) );
  NOR2_X1 U541 ( .A1(n758), .A2(n585), .ZN(n421) );
  NAND2_X1 U542 ( .A1(n424), .A2(n423), .ZN(n431) );
  NAND2_X1 U543 ( .A1(n432), .A2(n357), .ZN(n423) );
  OR2_X1 U544 ( .A1(n594), .A2(n595), .ZN(n426) );
  NAND2_X1 U545 ( .A1(n758), .A2(n585), .ZN(n427) );
  NAND2_X1 U546 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U547 ( .A1(n756), .A2(n585), .ZN(n429) );
  XNOR2_X1 U548 ( .A(n436), .B(n435), .ZN(n434) );
  INV_X1 U549 ( .A(KEYINPUT109), .ZN(n435) );
  NOR2_X1 U550 ( .A1(n690), .A2(n437), .ZN(n610) );
  NOR2_X1 U551 ( .A1(n673), .A2(n680), .ZN(n559) );
  XNOR2_X1 U552 ( .A(n496), .B(n440), .ZN(n568) );
  NAND2_X1 U553 ( .A1(n626), .A2(n730), .ZN(n666) );
  NAND2_X1 U554 ( .A1(n451), .A2(n730), .ZN(n450) );
  XNOR2_X2 U555 ( .A(n489), .B(KEYINPUT4), .ZN(n743) );
  XNOR2_X2 U556 ( .A(n459), .B(n458), .ZN(n489) );
  INV_X1 U557 ( .A(n683), .ZN(n447) );
  NAND2_X1 U558 ( .A1(n449), .A2(n354), .ZN(n571) );
  NAND2_X1 U559 ( .A1(n578), .A2(n670), .ZN(n551) );
  XNOR2_X2 U560 ( .A(n549), .B(n356), .ZN(n578) );
  NAND2_X1 U561 ( .A1(n450), .A2(n617), .ZN(n665) );
  OR2_X1 U562 ( .A1(n625), .A2(n606), .ZN(n748) );
  NOR2_X1 U563 ( .A1(n625), .A2(n452), .ZN(n451) );
  INV_X1 U564 ( .A(n606), .ZN(n453) );
  NAND2_X1 U565 ( .A1(n613), .A2(n563), .ZN(n455) );
  XOR2_X1 U566 ( .A(n479), .B(n478), .Z(n456) );
  XOR2_X1 U567 ( .A(G472), .B(KEYINPUT73), .Z(n457) );
  INV_X1 U568 ( .A(KEYINPUT74), .ZN(n595) );
  XNOR2_X1 U569 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n581) );
  XNOR2_X1 U570 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U571 ( .A(KEYINPUT48), .ZN(n602) );
  XNOR2_X1 U572 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U573 ( .A(n603), .B(n602), .ZN(n625) );
  BUF_X1 U574 ( .A(n489), .Z(n493) );
  BUF_X1 U575 ( .A(n669), .Z(n702) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n516) );
  INV_X1 U577 ( .A(KEYINPUT111), .ZN(n584) );
  XNOR2_X2 U578 ( .A(KEYINPUT65), .B(G143), .ZN(n459) );
  XOR2_X1 U579 ( .A(G104), .B(G107), .Z(n461) );
  XNOR2_X1 U580 ( .A(n461), .B(n460), .ZN(n545) );
  XOR2_X1 U581 ( .A(n545), .B(n515), .Z(n463) );
  NAND2_X1 U582 ( .A1(G227), .A2(n735), .ZN(n462) );
  XNOR2_X1 U583 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U584 ( .A(G469), .ZN(n465) );
  XNOR2_X1 U585 ( .A(n467), .B(G125), .ZN(n540) );
  XOR2_X1 U586 ( .A(n514), .B(G104), .Z(n472) );
  INV_X1 U587 ( .A(n469), .ZN(n470) );
  XOR2_X1 U588 ( .A(G113), .B(n470), .Z(n471) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n474), .B(n473), .ZN(n477) );
  XOR2_X1 U591 ( .A(KEYINPUT77), .B(n475), .Z(n504) );
  NAND2_X1 U592 ( .A1(G214), .A2(n504), .ZN(n476) );
  XNOR2_X1 U593 ( .A(n477), .B(n476), .ZN(n480) );
  XOR2_X1 U594 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n479) );
  XNOR2_X1 U595 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n478) );
  NAND2_X1 U596 ( .A1(n632), .A2(n534), .ZN(n484) );
  XOR2_X1 U597 ( .A(KEYINPUT13), .B(G475), .Z(n483) );
  XNOR2_X1 U598 ( .A(n484), .B(n483), .ZN(n587) );
  XNOR2_X1 U599 ( .A(G116), .B(G134), .ZN(n485) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n495) );
  XOR2_X1 U601 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n488) );
  NAND2_X1 U602 ( .A1(G234), .A2(n735), .ZN(n487) );
  XNOR2_X1 U603 ( .A(n488), .B(n487), .ZN(n507) );
  NAND2_X1 U604 ( .A1(G217), .A2(n507), .ZN(n494) );
  XOR2_X1 U605 ( .A(KEYINPUT104), .B(KEYINPUT102), .Z(n491) );
  XNOR2_X1 U606 ( .A(KEYINPUT103), .B(KEYINPUT105), .ZN(n490) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n492) );
  NOR2_X1 U608 ( .A1(G902), .A2(n722), .ZN(n496) );
  INV_X1 U609 ( .A(n568), .ZN(n586) );
  NAND2_X1 U610 ( .A1(n587), .A2(n586), .ZN(n658) );
  XNOR2_X1 U611 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U612 ( .A(n547), .B(n503), .Z(n506) );
  NAND2_X1 U613 ( .A1(n504), .A2(G210), .ZN(n505) );
  NAND2_X1 U614 ( .A1(G221), .A2(n507), .ZN(n513) );
  XOR2_X1 U615 ( .A(KEYINPUT24), .B(G110), .Z(n509) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U617 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n510) );
  XNOR2_X1 U618 ( .A(n515), .B(n514), .ZN(n745) );
  XNOR2_X1 U619 ( .A(n516), .B(n745), .ZN(n726) );
  NOR2_X1 U620 ( .A1(n726), .A2(G902), .ZN(n522) );
  XOR2_X1 U621 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n519) );
  NAND2_X1 U622 ( .A1(G234), .A2(n627), .ZN(n517) );
  XNOR2_X1 U623 ( .A(KEYINPUT20), .B(n517), .ZN(n523) );
  NAND2_X1 U624 ( .A1(n523), .A2(G217), .ZN(n518) );
  XNOR2_X1 U625 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U626 ( .A(n520), .B(KEYINPUT96), .ZN(n521) );
  NAND2_X1 U627 ( .A1(G221), .A2(n523), .ZN(n524) );
  XNOR2_X1 U628 ( .A(n524), .B(KEYINPUT21), .ZN(n680) );
  NAND2_X1 U629 ( .A1(G234), .A2(G237), .ZN(n525) );
  XNOR2_X1 U630 ( .A(n525), .B(KEYINPUT14), .ZN(n668) );
  INV_X1 U631 ( .A(G952), .ZN(n635) );
  NAND2_X1 U632 ( .A1(n735), .A2(n635), .ZN(n527) );
  OR2_X1 U633 ( .A1(n735), .A2(G902), .ZN(n526) );
  AND2_X1 U634 ( .A1(n527), .A2(n526), .ZN(n528) );
  AND2_X1 U635 ( .A1(n668), .A2(n528), .ZN(n553) );
  NAND2_X1 U636 ( .A1(G953), .A2(G900), .ZN(n747) );
  NAND2_X1 U637 ( .A1(n553), .A2(n747), .ZN(n529) );
  NOR2_X1 U638 ( .A1(n680), .A2(n350), .ZN(n530) );
  NAND2_X1 U639 ( .A1(n681), .A2(n530), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n565), .A2(n575), .ZN(n531) );
  XNOR2_X1 U641 ( .A(n531), .B(KEYINPUT107), .ZN(n532) );
  NOR2_X1 U642 ( .A1(n658), .A2(n532), .ZN(n535) );
  NAND2_X1 U643 ( .A1(n534), .A2(n533), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n548), .A2(G214), .ZN(n670) );
  NAND2_X1 U645 ( .A1(n535), .A2(n670), .ZN(n597) );
  NOR2_X1 U646 ( .A1(n683), .A2(n597), .ZN(n536) );
  XNOR2_X1 U647 ( .A(n536), .B(KEYINPUT43), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n735), .A2(G224), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n537), .B(KEYINPUT93), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n539), .B(n538), .ZN(n541) );
  XNOR2_X1 U651 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U652 ( .A(KEYINPUT16), .ZN(n543) );
  XNOR2_X1 U653 ( .A(n543), .B(G122), .ZN(n544) );
  XNOR2_X1 U654 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U655 ( .A(n547), .B(n546), .ZN(n736) );
  OR2_X1 U656 ( .A1(n550), .A2(n578), .ZN(n621) );
  XNOR2_X1 U657 ( .A(n621), .B(G140), .ZN(G42) );
  NAND2_X1 U658 ( .A1(G953), .A2(G898), .ZN(n552) );
  AND2_X1 U659 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U660 ( .A(KEYINPUT91), .B(KEYINPUT0), .ZN(n555) );
  INV_X1 U661 ( .A(KEYINPUT106), .ZN(n558) );
  XNOR2_X1 U662 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U663 ( .A(KEYINPUT80), .B(n565), .Z(n562) );
  NAND2_X1 U664 ( .A1(n683), .A2(n681), .ZN(n561) );
  NOR2_X1 U665 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U666 ( .A(n614), .B(G119), .Z(G21) );
  INV_X1 U667 ( .A(n565), .ZN(n573) );
  INV_X1 U668 ( .A(KEYINPUT79), .ZN(n569) );
  XNOR2_X1 U669 ( .A(n569), .B(KEYINPUT35), .ZN(n570) );
  XNOR2_X1 U670 ( .A(G122), .B(KEYINPUT127), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n367), .B(n572), .ZN(G24) );
  NOR2_X1 U672 ( .A1(n573), .A2(n683), .ZN(n574) );
  XNOR2_X1 U673 ( .A(KEYINPUT28), .B(n351), .ZN(n577) );
  INV_X1 U674 ( .A(n576), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n671), .A2(n670), .ZN(n674) );
  INV_X1 U676 ( .A(n658), .ZN(n655) );
  NAND2_X1 U677 ( .A1(n580), .A2(n670), .ZN(n582) );
  XNOR2_X1 U678 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n585) );
  OR2_X1 U679 ( .A1(n587), .A2(n586), .ZN(n661) );
  AND2_X1 U680 ( .A1(n661), .A2(n658), .ZN(n675) );
  NAND2_X1 U681 ( .A1(KEYINPUT47), .A2(n675), .ZN(n588) );
  XNOR2_X1 U682 ( .A(KEYINPUT84), .B(n588), .ZN(n589) );
  XNOR2_X1 U683 ( .A(n591), .B(KEYINPUT47), .ZN(n593) );
  INV_X1 U684 ( .A(n591), .ZN(n656) );
  NAND2_X1 U685 ( .A1(n656), .A2(n675), .ZN(n592) );
  NAND2_X1 U686 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U687 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U688 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n598) );
  XNOR2_X1 U689 ( .A(n599), .B(n598), .ZN(n600) );
  INV_X1 U690 ( .A(n661), .ZN(n652) );
  NAND2_X1 U691 ( .A1(n604), .A2(n652), .ZN(n605) );
  XOR2_X1 U692 ( .A(KEYINPUT113), .B(n605), .Z(n755) );
  NAND2_X1 U693 ( .A1(n755), .A2(n621), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n690) );
  AND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n650) );
  INV_X1 U696 ( .A(KEYINPUT82), .ZN(n619) );
  INV_X1 U697 ( .A(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n755), .A2(KEYINPUT2), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n618), .A2(KEYINPUT82), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n619), .A2(n755), .ZN(n620) );
  AND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U704 ( .A(n627), .ZN(n628) );
  INV_X1 U705 ( .A(KEYINPUT66), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n716), .A2(G475), .ZN(n634) );
  XNOR2_X1 U707 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n636) );
  NOR2_X2 U710 ( .A1(n636), .A2(n729), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U712 ( .A1(n716), .A2(G472), .ZN(n640) );
  XOR2_X1 U713 ( .A(KEYINPUT62), .B(n638), .Z(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X2 U715 ( .A1(n641), .A2(n729), .ZN(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(G57) );
  NOR2_X1 U718 ( .A1(n658), .A2(n647), .ZN(n644) );
  XOR2_X1 U719 ( .A(G104), .B(n644), .Z(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n646) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT27), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n661), .A2(n647), .ZN(n648) );
  XOR2_X1 U724 ( .A(n649), .B(n648), .Z(G9) );
  XNOR2_X1 U725 ( .A(G110), .B(n650), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT115), .ZN(G12) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  NAND2_X1 U728 ( .A1(n656), .A2(n652), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(G30) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(G146), .ZN(G48) );
  NOR2_X1 U732 ( .A1(n658), .A2(n660), .ZN(n659) );
  XOR2_X1 U733 ( .A(G113), .B(n659), .Z(G15) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U735 ( .A(G116), .B(n662), .Z(G18) );
  XNOR2_X1 U736 ( .A(n355), .B(KEYINPUT37), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(KEYINPUT116), .ZN(n664) );
  XNOR2_X1 U738 ( .A(G125), .B(n664), .ZN(G27) );
  NAND2_X1 U739 ( .A1(n665), .A2(n348), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n667), .B(KEYINPUT85), .ZN(n706) );
  NAND2_X1 U741 ( .A1(G952), .A2(n668), .ZN(n699) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(n678), .Z(n679) );
  NAND2_X1 U747 ( .A1(n702), .A2(n679), .ZN(n696) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT49), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U753 ( .A(n689), .B(KEYINPUT118), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n693) );
  XNOR2_X1 U755 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n692) );
  XNOR2_X1 U756 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n701), .A2(n694), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U759 ( .A(KEYINPUT52), .B(n697), .Z(n698) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U761 ( .A(n700), .B(KEYINPUT121), .ZN(n704) );
  NAND2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n735), .A2(n707), .ZN(n708) );
  XOR2_X1 U766 ( .A(KEYINPUT53), .B(n708), .Z(G75) );
  AND2_X2 U767 ( .A1(n716), .A2(G210), .ZN(n713) );
  XOR2_X1 U768 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n710) );
  XOR2_X1 U769 ( .A(n710), .B(KEYINPUT55), .Z(n711) );
  XOR2_X1 U770 ( .A(n709), .B(n711), .Z(n712) );
  XNOR2_X1 U771 ( .A(KEYINPUT56), .B(n715), .ZN(G51) );
  NAND2_X1 U772 ( .A1(n725), .A2(G469), .ZN(n720) );
  XOR2_X1 U773 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  XNOR2_X1 U774 ( .A(n717), .B(KEYINPUT123), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n729), .A2(n721), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n725), .A2(G478), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n729), .A2(n724), .ZN(G63) );
  NAND2_X1 U779 ( .A1(n725), .A2(G217), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(G66) );
  NAND2_X1 U782 ( .A1(n730), .A2(n735), .ZN(n734) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n741) );
  NOR2_X1 U787 ( .A1(G898), .A2(n735), .ZN(n738) );
  XOR2_X1 U788 ( .A(n736), .B(G101), .Z(n737) );
  NOR2_X1 U789 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U790 ( .A(KEYINPUT125), .B(n739), .Z(n740) );
  XNOR2_X1 U791 ( .A(n741), .B(n740), .ZN(G69) );
  XOR2_X1 U792 ( .A(n743), .B(n742), .Z(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n749) );
  XNOR2_X1 U794 ( .A(n749), .B(G227), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n752) );
  XOR2_X1 U796 ( .A(n749), .B(n748), .Z(n750) );
  NOR2_X1 U797 ( .A1(G953), .A2(n750), .ZN(n751) );
  NOR2_X1 U798 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U799 ( .A(n753), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U800 ( .A(G134), .B(KEYINPUT117), .Z(n754) );
  XNOR2_X1 U801 ( .A(n755), .B(n754), .ZN(G36) );
  XOR2_X1 U802 ( .A(n756), .B(G137), .Z(G39) );
  XNOR2_X1 U803 ( .A(n757), .B(G143), .ZN(G45) );
  XOR2_X1 U804 ( .A(n758), .B(G131), .Z(G33) );
endmodule

