//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(KEYINPUT64), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT64), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n190), .A3(new_n192), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n193), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n190), .A2(new_n192), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G224), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n203), .B(new_n209), .C1(new_n211), .C2(G953), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(G110), .B(G122), .Z(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT76), .B(G101), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n225), .A3(new_n221), .A4(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n221), .A2(G104), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n224), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n223), .A2(new_n226), .A3(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(G101), .A3(new_n230), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n219), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(G113), .C1(KEYINPUT5), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n217), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n241), .A2(new_n218), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G107), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n245), .B2(new_n227), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n229), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n216), .B1(new_n236), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT6), .ZN(new_n250));
  INV_X1    g064(.A(new_n219), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n229), .A2(new_n230), .B1(new_n232), .B2(G101), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n232), .A2(G101), .A3(new_n230), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n216), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n229), .A2(new_n246), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n242), .A3(new_n240), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT81), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n254), .B2(new_n257), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT6), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT82), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n236), .A2(new_n248), .A3(new_n216), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n264), .B2(new_n260), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n249), .B2(KEYINPUT81), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n215), .B(new_n250), .C1(new_n263), .C2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n216), .B(KEYINPUT8), .Z(new_n271));
  AOI21_X1  g085(.A(KEYINPUT83), .B1(new_n243), .B2(new_n247), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n248), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n243), .A2(KEYINPUT83), .A3(new_n247), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n213), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n258), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n188), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n215), .ZN(new_n282));
  INV_X1    g096(.A(new_n250), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT82), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n268), .B1(new_n265), .B2(new_n267), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n280), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n187), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G214), .B1(G237), .B2(G902), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n290), .B(KEYINPUT80), .Z(new_n291));
  AND2_X1   g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n234), .A2(new_n235), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT10), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n197), .B2(new_n200), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n296), .A2(new_n208), .B1(new_n256), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(G143), .B2(new_n189), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n198), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n193), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n200), .B(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n247), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n310), .A2(KEYINPUT79), .A3(KEYINPUT10), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n303), .A2(new_n305), .B1(new_n190), .B2(new_n192), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n200), .B(KEYINPUT77), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n256), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(new_n297), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n299), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G137), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT11), .A3(G134), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G131), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n320), .A2(new_n322), .A3(new_n326), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n325), .A2(KEYINPUT66), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n317), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  INV_X1    g149(.A(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n335), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n208), .B1(new_n252), .B2(new_n253), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n298), .A2(new_n256), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n315), .A2(new_n312), .A3(new_n297), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT79), .B1(new_n310), .B2(KEYINPUT10), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n339), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n332), .B(new_n299), .C1(new_n311), .C2(new_n316), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n247), .A2(new_n200), .A3(new_n197), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT12), .B(new_n328), .C1(new_n349), .C2(new_n310), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n332), .B1(new_n315), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n338), .B(KEYINPUT73), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n334), .A2(new_n346), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G469), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(G469), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n338), .B1(new_n334), .B2(new_n347), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n347), .A2(new_n338), .A3(new_n352), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n357), .B(new_n279), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n295), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  AND4_X1   g176(.A1(G143), .A2(new_n362), .A3(new_n336), .A4(G214), .ZN(new_n363));
  NOR2_X1   g177(.A1(G237), .A2(G953), .ZN(new_n364));
  AOI21_X1  g178(.A(G143), .B1(new_n364), .B2(G214), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT18), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n326), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n336), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n191), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n364), .A2(G143), .A3(G214), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(new_n372), .C1(new_n368), .C2(new_n326), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT84), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n202), .A2(G140), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n189), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n202), .A2(G140), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n375), .B2(G125), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n202), .A2(KEYINPUT69), .A3(G140), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n383), .B2(new_n189), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n371), .A2(new_n372), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT18), .A3(G131), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n369), .A2(new_n374), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n363), .B2(new_n365), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n371), .A2(new_n326), .A3(new_n372), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT19), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n376), .A2(new_n377), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n189), .B(new_n392), .C1(new_n383), .C2(new_n391), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n379), .A2(KEYINPUT16), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n202), .A2(KEYINPUT69), .A3(G140), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT69), .B1(new_n202), .B2(G140), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n376), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n390), .B(new_n393), .C1(new_n398), .C2(new_n189), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n387), .A2(KEYINPUT85), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n387), .B2(new_n399), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n244), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT86), .B1(new_n388), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n385), .A2(new_n407), .A3(KEYINPUT17), .A4(G131), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(new_n408), .C1(KEYINPUT17), .C2(new_n390), .ZN(new_n409));
  INV_X1    g223(.A(new_n394), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n383), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G146), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n410), .B(new_n189), .C1(new_n383), .C2(new_n411), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n403), .B(new_n387), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT87), .B1(new_n404), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n404), .B2(new_n417), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI221_X1 g236(.A(new_n419), .B1(KEYINPUT87), .B2(KEYINPUT20), .C1(new_n404), .C2(new_n417), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n409), .A2(new_n415), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n403), .B1(new_n425), .B2(new_n387), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n279), .B1(new_n426), .B2(new_n417), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G475), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n293), .A2(new_n429), .A3(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n198), .A2(G143), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n319), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n191), .A2(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n432), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n436), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G116), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G122), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(new_n440), .A3(G122), .ZN(new_n443));
  INV_X1    g257(.A(G122), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT88), .B1(new_n444), .B2(G116), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n221), .B(new_n441), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n432), .A3(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n436), .A2(new_n319), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n443), .A2(new_n445), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n444), .B2(G116), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT89), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(KEYINPUT89), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n452), .B1(new_n458), .B2(G107), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n431), .B1(new_n449), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n454), .B1(new_n443), .B2(new_n445), .ZN(new_n462));
  OAI21_X1  g276(.A(G107), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n451), .A2(new_n450), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n446), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n448), .A2(new_n446), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n438), .A3(new_n437), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(new_n430), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n468), .A3(KEYINPUT90), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n467), .A3(new_n470), .A4(new_n430), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n471), .A3(new_n279), .ZN(new_n472));
  INV_X1    g286(.A(G478), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n469), .A2(new_n471), .A3(new_n279), .A4(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n428), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT92), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n279), .B(new_n336), .C1(G234), .C2(G237), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n336), .A2(G952), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G234), .B2(G237), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n424), .A2(new_n482), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n292), .A2(new_n361), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G472), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n330), .A2(new_n208), .A3(new_n331), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n319), .A2(G137), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n321), .A2(G134), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n327), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n197), .B2(new_n200), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n219), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n495), .A2(KEYINPUT28), .A3(new_n219), .A4(new_n501), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n364), .A2(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G101), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n495), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n251), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n506), .A2(KEYINPUT29), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n279), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n325), .A2(new_n327), .B1(new_n205), .B2(new_n207), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n500), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT65), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n495), .A2(KEYINPUT30), .A3(new_n501), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(new_n515), .C1(new_n500), .C2(new_n516), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n518), .A2(new_n519), .A3(new_n251), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n502), .ZN(new_n523));
  INV_X1    g337(.A(new_n510), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n251), .B1(new_n500), .B2(new_n516), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n504), .A2(new_n527), .A3(new_n505), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n525), .B(new_n526), .C1(new_n524), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n494), .B1(new_n514), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n502), .A3(new_n510), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n524), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n522), .A2(new_n534), .A3(new_n502), .A4(new_n510), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n494), .A3(new_n279), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(KEYINPUT32), .A3(new_n494), .A4(new_n279), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(KEYINPUT67), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n537), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT32), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n530), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n238), .A2(G128), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT68), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT68), .B1(new_n238), .B2(G128), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n198), .A2(G119), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  OAI22_X1  g370(.A1(new_n553), .A2(G110), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n413), .A2(new_n557), .A3(new_n378), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(G110), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n413), .B2(new_n414), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT70), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n415), .A2(new_n561), .A3(new_n560), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n558), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT22), .B(G137), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n336), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n558), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n279), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n573), .A2(new_n279), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n429), .B1(G234), .B2(new_n279), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G902), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT72), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n573), .ZN(new_n586));
  INV_X1    g400(.A(new_n574), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n581), .A2(new_n582), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n545), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n493), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(new_n224), .Z(G3));
  NOR2_X1   g407(.A1(new_n590), .A2(new_n295), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n356), .A2(new_n360), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n536), .A2(new_n279), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n494), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n290), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n281), .B2(new_n288), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n422), .A2(new_n423), .A3(new_n428), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n469), .A2(new_n471), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n460), .A2(new_n468), .A3(KEYINPUT33), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n279), .A4(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n472), .A2(KEYINPUT93), .A3(new_n473), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT93), .B1(new_n472), .B2(new_n473), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n487), .B2(new_n490), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  NAND2_X1  g428(.A1(new_n479), .A2(new_n481), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n420), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n401), .A2(new_n403), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n416), .B1(new_n619), .B2(new_n400), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n419), .A3(new_n616), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n615), .A2(new_n428), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n491), .B(KEYINPUT95), .Z(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n601), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G107), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n571), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT97), .Z(new_n631));
  AND3_X1   g445(.A1(new_n564), .A2(new_n567), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n564), .B2(new_n567), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n585), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(new_n585), .C1(new_n632), .C2(new_n633), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n581), .B2(new_n582), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n493), .A2(new_n597), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT37), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G12));
  NAND2_X1  g458(.A1(new_n541), .A2(new_n544), .ZN(new_n645));
  INV_X1    g459(.A(new_n530), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n640), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n489), .B1(new_n486), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n622), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n250), .B1(new_n263), .B2(new_n269), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n188), .B(new_n280), .C1(new_n652), .C2(new_n282), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n187), .B1(new_n286), .B2(new_n287), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n290), .B(new_n651), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n289), .A2(new_n657), .A3(new_n290), .A4(new_n651), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n656), .A2(new_n658), .A3(new_n361), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n198), .ZN(G30));
  INV_X1    g475(.A(new_n531), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n510), .B1(new_n512), .B2(new_n502), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n279), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G472), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n645), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n289), .B(KEYINPUT38), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n650), .B(KEYINPUT39), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n361), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n640), .A2(new_n599), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n602), .A2(new_n615), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OR4_X1    g491(.A1(new_n667), .A2(new_n669), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n650), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n602), .A2(new_n609), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n361), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n290), .B1(new_n653), .B2(new_n654), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n647), .A2(new_n640), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  OAI21_X1  g500(.A(new_n279), .B1(new_n358), .B2(new_n359), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n294), .A3(new_n360), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n600), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n545), .A2(new_n690), .A3(new_n590), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n611), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n624), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n545), .A2(new_n639), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n600), .A2(new_n492), .A3(new_n689), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n697), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT101), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n238), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(new_n623), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n506), .A2(new_n512), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n524), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n532), .A3(new_n535), .ZN(new_n707));
  NOR2_X1   g521(.A1(G472), .A2(G902), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n596), .A2(G472), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n689), .A2(new_n589), .A3(new_n704), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n289), .A2(new_n711), .A3(new_n290), .A4(new_n676), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n676), .B(new_n290), .C1(new_n653), .C2(new_n654), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n703), .B(new_n710), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n712), .ZN(new_n716));
  INV_X1    g530(.A(new_n710), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT103), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n444), .ZN(G24));
  INV_X1    g534(.A(new_n689), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n683), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n640), .A2(new_n709), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n681), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NOR2_X1   g539(.A1(new_n289), .A2(new_n599), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n361), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n681), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(KEYINPUT42), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n591), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n361), .A3(new_n681), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n646), .A2(new_n539), .A3(new_n540), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n589), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT42), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n326), .ZN(G33));
  NAND3_X1  g551(.A1(new_n728), .A2(new_n591), .A3(new_n651), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  OR2_X1    g553(.A1(new_n355), .A2(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n355), .A2(KEYINPUT45), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(G469), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(G469), .A2(G902), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n360), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n294), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n609), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n602), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n602), .B2(KEYINPUT104), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n751), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n597), .A2(new_n639), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n726), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n754), .A2(KEYINPUT44), .A3(new_n755), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n749), .A2(new_n671), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  OR2_X1    g575(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT106), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n647), .A2(new_n757), .A3(new_n589), .A4(new_n729), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  AND2_X1   g583(.A1(new_n688), .A2(new_n360), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT49), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n594), .A2(new_n291), .A3(new_n751), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(KEYINPUT107), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n667), .A4(new_n669), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n726), .A2(new_n689), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT115), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n589), .A3(new_n489), .A4(new_n667), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT116), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n602), .A3(new_n609), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n754), .A2(new_n489), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n734), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT48), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n589), .A2(new_n709), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n488), .B1(new_n789), .B2(new_n722), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n780), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT118), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n764), .A2(new_n766), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n770), .A2(new_n295), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT114), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n757), .B(new_n788), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n779), .A2(new_n424), .A3(new_n428), .A4(new_n750), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n668), .A2(new_n290), .A3(new_n721), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n789), .A2(KEYINPUT50), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  INV_X1    g614(.A(new_n798), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n788), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n799), .A2(new_n802), .B1(new_n782), .B2(new_n723), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n796), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n793), .A2(new_n806), .A3(new_n794), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n726), .A3(new_n789), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n793), .B2(new_n794), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n811));
  OAI221_X1 g625(.A(new_n792), .B1(new_n805), .B2(KEYINPUT51), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n482), .A2(new_n621), .A3(new_n618), .A4(new_n680), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT108), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n697), .A2(new_n814), .B1(new_n681), .B2(new_n723), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n738), .B1(new_n815), .B2(new_n727), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(KEYINPUT109), .B(new_n738), .C1(new_n815), .C2(new_n727), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n650), .B(KEYINPUT110), .Z(new_n822));
  NAND3_X1  g636(.A1(new_n361), .A2(new_n639), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n645), .B2(new_n665), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n716), .A2(KEYINPUT111), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT111), .B1(new_n716), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n685), .B(new_n724), .C1(new_n648), .C2(new_n659), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n716), .A2(new_n824), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n716), .A2(new_n824), .A3(KEYINPUT111), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n828), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n615), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n610), .B1(new_n838), .B2(new_n602), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n598), .A2(new_n292), .A3(new_n704), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n641), .A3(new_n592), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(KEYINPUT112), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n820), .A2(new_n837), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n692), .B(new_n695), .C1(new_n715), .C2(new_n718), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n701), .A3(new_n736), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n837), .A2(new_n820), .A3(new_n842), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n843), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n841), .B1(new_n829), .B2(new_n836), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n820), .A4(new_n847), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n845), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n837), .A2(new_n820), .A3(new_n842), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n853), .A2(KEYINPUT112), .A3(new_n843), .A4(new_n847), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n852), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT113), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n845), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  INV_X1    g676(.A(new_n854), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n857), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n812), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n775), .B1(new_n867), .B2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n336), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g685(.A(G902), .B1(new_n852), .B2(new_n854), .ZN(new_n872));
  INV_X1    g686(.A(G210), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n652), .B(new_n282), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n188), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n870), .B(new_n877), .C1(new_n881), .C2(new_n882), .ZN(G51));
  INV_X1    g697(.A(new_n742), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n743), .B(KEYINPUT57), .Z(new_n886));
  AOI21_X1  g700(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n855), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n358), .B2(new_n359), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n870), .B1(new_n885), .B2(new_n889), .ZN(G54));
  NAND2_X1  g704(.A1(KEYINPUT58), .A2(G475), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n878), .B2(new_n879), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n620), .ZN(new_n893));
  INV_X1    g707(.A(new_n870), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n892), .B2(new_n620), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n859), .A2(new_n866), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n604), .A2(new_n605), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n898), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n852), .B2(new_n854), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n864), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n894), .B1(new_n907), .B2(KEYINPUT120), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n909), .B(new_n905), .C1(new_n864), .C2(new_n906), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n903), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n904), .B1(new_n887), .B2(new_n855), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT121), .A4(new_n894), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n902), .B1(new_n911), .B2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(new_n861), .A2(new_n863), .ZN(new_n917));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  AOI21_X1  g733(.A(new_n588), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n919), .B1(new_n632), .B2(new_n633), .C1(new_n852), .C2(new_n854), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n894), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n920), .A2(new_n922), .B1(KEYINPUT122), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(KEYINPUT122), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G66));
  AOI21_X1  g740(.A(new_n336), .B1(new_n484), .B2(G224), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n846), .A2(new_n841), .A3(new_n701), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n336), .ZN(new_n929));
  INV_X1    g743(.A(G898), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n652), .B1(new_n930), .B2(G953), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  AOI21_X1  g746(.A(new_n336), .B1(G227), .B2(G900), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n649), .A2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n749), .A2(new_n671), .A3(new_n783), .ZN(new_n937));
  INV_X1    g751(.A(new_n716), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n738), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n736), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n768), .A2(new_n940), .A3(new_n760), .A4(new_n835), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n936), .B1(new_n941), .B2(new_n336), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(KEYINPUT125), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n392), .B1(new_n383), .B2(new_n391), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n942), .B2(KEYINPUT125), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  INV_X1    g763(.A(new_n672), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n591), .A2(new_n839), .A3(new_n950), .A4(new_n726), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n768), .A2(new_n760), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n678), .A2(new_n835), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n336), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n946), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n933), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n957), .B(new_n933), .C1(new_n943), .C2(new_n947), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT126), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n941), .B2(new_n928), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n523), .B(KEYINPUT127), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n510), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n870), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n952), .A2(new_n928), .A3(new_n954), .ZN(new_n969));
  INV_X1    g783(.A(new_n964), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n966), .A2(new_n510), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n525), .A2(new_n531), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n963), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n856), .B2(new_n975), .ZN(G57));
endmodule


