//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n467), .B2(new_n474), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n467), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n482), .A2(G124), .B1(G136), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT68), .Z(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n463), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G102), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n474), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n479), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n503), .B(new_n505), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT69), .B(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n509), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  AND3_X1   g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT70), .B(G51), .Z(new_n523));
  OAI221_X1 g098(.A(new_n521), .B1(KEYINPUT7), .B2(new_n522), .C1(new_n513), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n506), .A2(G63), .ZN(new_n525));
  NAND3_X1  g100(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n508), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n513), .A2(new_n531), .B1(new_n532), .B2(new_n515), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n513), .A2(new_n537), .B1(new_n538), .B2(new_n515), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT71), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n541), .B1(new_n538), .B2(new_n515), .C1(new_n513), .C2(new_n537), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n536), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G860), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT72), .Z(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n520), .A2(G91), .ZN(new_n553));
  OAI211_X1 g128(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OAI221_X1 g132(.A(new_n553), .B1(new_n556), .B2(KEYINPUT9), .C1(new_n557), .C2(new_n508), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n554), .A2(new_n555), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n559), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n558), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  OR2_X1    g138(.A1(new_n506), .A2(G74), .ZN(new_n564));
  INV_X1    g139(.A(new_n513), .ZN(new_n565));
  AOI22_X1  g140(.A1(G651), .A2(new_n564), .B1(new_n565), .B2(G49), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n515), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n520), .A2(KEYINPUT74), .A3(G87), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n506), .A2(G61), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n508), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g149(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n515), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT75), .ZN(G305));
  AOI22_X1  g154(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n508), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n513), .A2(new_n582), .B1(new_n583), .B2(new_n515), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n503), .A2(new_n505), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n565), .A2(G54), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT10), .B1(new_n515), .B2(new_n592), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G321));
  NAND2_X1  g174(.A1(G299), .A2(new_n596), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g177(.A(new_n595), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g181(.A1(new_n544), .A2(new_n596), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n595), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n596), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g185(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT78), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n479), .A2(new_n494), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n612), .B(new_n613), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n482), .A2(G123), .B1(G135), .B2(new_n483), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT80), .Z(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n635), .B(new_n638), .Z(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(G14), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n643), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT18), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  AOI22_X1  g237(.A1(new_n660), .A2(new_n661), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n657), .A2(new_n662), .A3(new_n659), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n663), .B(new_n664), .C1(new_n661), .C2(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1981), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT85), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  NOR2_X1   g247(.A1(G25), .A2(G29), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n482), .A2(G119), .B1(G131), .B2(new_n483), .ZN(new_n674));
  OR2_X1    g249(.A1(G95), .A2(G2105), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n673), .B1(new_n678), .B2(G29), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT35), .B(G1991), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G24), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n585), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1986), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT32), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G1971), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(G1971), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n694), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n689), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n686), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT36), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n621), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT89), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n706), .B1(new_n715), .B2(G34), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(G34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n476), .B2(new_n706), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G5), .B2(G16), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n725), .A2(G5), .A3(G16), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n726), .B(new_n727), .C1(G301), .C2(new_n695), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n603), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G4), .B2(G16), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n724), .B(new_n730), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G19), .B(new_n544), .S(G16), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G1341), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT31), .B(G11), .Z(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n738), .A2(G28), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(G28), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n739), .A2(new_n740), .A3(G29), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G21), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G168), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n737), .B(new_n741), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n714), .A2(new_n734), .A3(new_n736), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n728), .A2(new_n729), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n735), .A2(G1341), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT26), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n482), .B2(G129), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n494), .A2(G105), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n483), .A2(G141), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  OAI22_X1  g335(.A1(new_n712), .A2(new_n713), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n706), .A2(G33), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G103), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n483), .A2(G139), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n764), .B(new_n765), .C1(new_n474), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT87), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(new_n706), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n695), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT93), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n706), .A2(G26), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n482), .A2(G128), .B1(G140), .B2(new_n483), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n777), .B1(new_n782), .B2(new_n706), .ZN(new_n783));
  MUX2_X1   g358(.A(new_n777), .B(new_n783), .S(KEYINPUT28), .Z(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n759), .A2(new_n760), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n706), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n706), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n771), .A2(new_n776), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n761), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n705), .A2(new_n708), .A3(new_n750), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n744), .A2(new_n745), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n733), .A2(new_n731), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(G311));
  NAND2_X1  g374(.A1(new_n750), .A2(new_n795), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n704), .A2(KEYINPUT36), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n704), .A2(KEYINPUT36), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n797), .ZN(new_n804));
  INV_X1    g379(.A(new_n798), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n708), .ZN(G150));
  AOI22_X1  g381(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n508), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n513), .A2(new_n809), .B1(new_n810), .B2(new_n515), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n808), .B2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n545), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n816), .A2(new_n544), .ZN(new_n821));
  INV_X1    g396(.A(new_n812), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(new_n536), .C1(new_n540), .C2(new_n543), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT95), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n816), .A2(new_n544), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n595), .A2(new_n604), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n829), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n820), .B1(new_n833), .B2(G860), .ZN(G145));
  NAND2_X1  g409(.A1(new_n482), .A2(G130), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n483), .A2(G142), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT98), .Z(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n614), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n677), .B(KEYINPUT100), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT101), .ZN(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n757), .B(new_n781), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(G164), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(G164), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n769), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n767), .A3(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n846), .A2(new_n850), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n621), .B(new_n476), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n488), .B(new_n863), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n848), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n860), .A3(new_n864), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  NAND2_X1  g449(.A1(G299), .A2(new_n603), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n558), .A2(new_n560), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n595), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(KEYINPUT103), .A3(new_n877), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n876), .A2(KEYINPUT103), .A3(new_n595), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n877), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n825), .A2(new_n608), .A3(new_n828), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n608), .B1(new_n825), .B2(new_n828), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n881), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n880), .B(KEYINPUT104), .ZN(new_n889));
  INV_X1    g464(.A(new_n887), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G305), .B(G303), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(new_n585), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(new_n891), .A3(new_n874), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n896), .ZN(new_n899));
  INV_X1    g474(.A(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G868), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n816), .A2(G868), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n873), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n596), .B1(new_n898), .B2(new_n901), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n907), .A2(KEYINPUT105), .A3(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(G295));
  NAND2_X1  g484(.A1(new_n903), .A2(new_n905), .ZN(G331));
  XNOR2_X1  g485(.A(G168), .B(G171), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n828), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n827), .B1(new_n826), .B2(new_n823), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n825), .A2(new_n828), .A3(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n880), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n884), .B1(new_n919), .B2(new_n883), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n825), .A2(KEYINPUT106), .A3(new_n828), .A4(new_n911), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n825), .A2(new_n925), .A3(new_n828), .A4(new_n911), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n880), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n896), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n924), .A2(new_n926), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n899), .B(new_n922), .C1(new_n929), .C2(new_n880), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n880), .A2(new_n883), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n926), .A2(new_n924), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n889), .B1(new_n918), .B2(new_n921), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n896), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n931), .A4(new_n930), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n933), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n930), .A2(new_n931), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n932), .A2(new_n939), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT44), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(G397));
  AND2_X1   g524(.A1(new_n498), .A2(new_n499), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n494), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n470), .A2(new_n475), .A3(G40), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n757), .B(G1996), .Z(new_n956));
  XNOR2_X1  g531(.A(new_n781), .B(new_n785), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n677), .A2(new_n681), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n782), .A2(new_n785), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n955), .A2(G1996), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT46), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n955), .B1(new_n957), .B2(new_n758), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n956), .A2(new_n957), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n677), .A2(new_n681), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n967), .A2(new_n958), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n955), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  NOR2_X1   g548(.A1(G290), .A2(G1986), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT48), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n961), .B(new_n966), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n954), .B1(new_n952), .B2(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n479), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n495), .B1(new_n980), .B2(new_n474), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n498), .A2(new_n499), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT45), .B(new_n979), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n745), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT50), .B(new_n979), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT50), .B1(new_n500), .B2(new_n979), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n723), .B(new_n954), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(G168), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(KEYINPUT51), .A3(G8), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(KEYINPUT121), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n985), .A2(new_n989), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(G8), .A3(G286), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(KEYINPUT120), .A3(G8), .A4(G286), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n991), .A2(new_n1002), .A3(new_n992), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n995), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n995), .A2(new_n1001), .A3(new_n1006), .A4(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n470), .A2(new_n475), .A3(G40), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n952), .A2(new_n1015), .A3(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n983), .A2(KEYINPUT109), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1010), .B1(new_n1018), .B2(G2078), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n954), .B1(new_n987), .B2(new_n988), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n729), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1010), .A2(G2078), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n983), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G171), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT55), .Z(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1018), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1012), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1011), .B1(new_n1031), .B2(new_n986), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT111), .B(G2090), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1027), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n578), .B2(new_n1038), .ZN(new_n1039));
  NOR4_X1   g614(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT112), .A4(G1981), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1039), .A2(new_n1040), .B1(new_n1038), .B2(new_n578), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n952), .A2(new_n954), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  OAI221_X1 g620(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n578), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1048), .B2(G288), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1045), .B(new_n1051), .C1(new_n1048), .C2(G288), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1036), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1018), .A2(new_n1056), .A3(new_n1028), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1034), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(G8), .A3(new_n1027), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1054), .A2(KEYINPUT123), .A3(new_n1059), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1025), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1005), .A2(new_n1065), .A3(new_n1007), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1009), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1047), .A2(new_n1048), .A3(new_n691), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1045), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1059), .B2(new_n1053), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1027), .B1(new_n1058), .B2(G8), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1072), .A2(KEYINPUT113), .A3(new_n1053), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT113), .B1(new_n1072), .B2(new_n1053), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n996), .A2(G8), .A3(G168), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1073), .A2(new_n1059), .A3(new_n1074), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1060), .B2(new_n1076), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1067), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1022), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1019), .A2(new_n1021), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n1086), .B2(new_n1025), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(G171), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1019), .A2(G301), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(KEYINPUT54), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1089), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1008), .A2(new_n1083), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1008), .A2(new_n1083), .A3(KEYINPUT125), .A4(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  NAND3_X1  g675(.A1(G299), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n876), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT116), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT114), .B(G1956), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1020), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1106), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1020), .A2(new_n731), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1044), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n785), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n595), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1112), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1111), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1105), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1122), .A2(new_n1113), .A3(new_n1125), .A4(KEYINPUT61), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1121), .A2(new_n1105), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1112), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1116), .B1(new_n1032), .B2(G1348), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n603), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1117), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1131), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1018), .A2(G1996), .B1(new_n1115), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n540), .A2(new_n543), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(KEYINPUT117), .A3(new_n536), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT59), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1130), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1100), .B(new_n1118), .C1(new_n1127), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1135), .B1(new_n1145), .B2(new_n1128), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n1124), .A3(new_n1141), .A4(new_n1126), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1100), .B1(new_n1147), .B2(new_n1118), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1082), .B1(new_n1099), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n970), .B1(G1986), .B2(G290), .ZN(new_n1151));
  INV_X1    g726(.A(new_n974), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n955), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n977), .B1(new_n1150), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g729(.A(new_n460), .B1(new_n866), .B2(new_n870), .ZN(new_n1156));
  NOR3_X1   g730(.A1(G401), .A2(G227), .A3(G229), .ZN(new_n1157));
  NAND4_X1  g731(.A1(new_n1156), .A2(new_n941), .A3(new_n942), .A4(new_n1157), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


