//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G110), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT24), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n196), .B2(new_n198), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n188), .B2(G119), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(KEYINPUT75), .A3(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR4_X1    g019(.A1(new_n194), .A2(new_n200), .A3(new_n201), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT16), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n212), .A3(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT66), .B(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT23), .B1(new_n188), .B2(G119), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n193), .B2(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n223), .B2(G110), .ZN(new_n224));
  AOI211_X1 g038(.A(KEYINPUT77), .B(new_n195), .C1(new_n220), .C2(new_n222), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n206), .B(new_n217), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n194), .A2(new_n205), .B1(new_n200), .B2(new_n201), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(G110), .B2(new_n223), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT78), .A4(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(G125), .B(G140), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n214), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(new_n230), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G137), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n236), .B(new_n238), .Z(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n226), .A2(new_n234), .A3(KEYINPUT79), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n239), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n187), .B1(new_n247), .B2(G902), .ZN(new_n248));
  INV_X1    g062(.A(new_n244), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT79), .B1(new_n226), .B2(new_n234), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n240), .ZN(new_n252));
  INV_X1    g066(.A(G902), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G217), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(G234), .B2(new_n253), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G902), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n255), .A2(new_n257), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT32), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n214), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(G143), .B2(new_n214), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n219), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND4_X1   g086(.A1(new_n269), .A2(new_n271), .A3(new_n262), .A4(new_n264), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(G137), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n277), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n276), .A2(G137), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n278), .A2(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(G131), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n285), .A3(KEYINPUT64), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n274), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n262), .A2(new_n264), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT0), .B(G128), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n270), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G131), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n282), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n261), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n193), .A2(G116), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(G119), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n193), .A2(KEYINPUT67), .A3(G116), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G113), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n301), .A2(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT67), .B1(new_n193), .B2(G116), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n301), .A3(G119), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n286), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n296), .A2(new_n282), .ZN(new_n319));
  INV_X1    g133(.A(new_n294), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n274), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT68), .B1(new_n321), .B2(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n271), .A2(new_n262), .A3(new_n264), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n270), .A2(new_n269), .A3(new_n271), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n286), .B1(new_n326), .B2(new_n268), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  NOR4_X1   g142(.A1(new_n327), .A2(new_n297), .A3(new_n328), .A4(new_n261), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n298), .B(new_n317), .C1(new_n322), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  INV_X1    g145(.A(new_n317), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  NOR2_X1   g148(.A1(G237), .A2(G953), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G210), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n331), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n317), .B1(new_n290), .B2(new_n297), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n321), .A2(KEYINPUT28), .A3(new_n332), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n339), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n274), .A2(new_n288), .A3(new_n289), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n319), .A2(new_n320), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT30), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n192), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n324), .A2(new_n325), .B1(new_n355), .B2(new_n265), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n352), .B(KEYINPUT30), .C1(new_n286), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n328), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n321), .A2(KEYINPUT68), .A3(KEYINPUT30), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n340), .B1(new_n360), .B2(new_n317), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT70), .B1(new_n361), .B2(new_n331), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n331), .B1(new_n330), .B2(new_n341), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n350), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT71), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n260), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n361), .A2(new_n331), .B1(new_n348), .B2(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n330), .A2(new_n341), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n364), .B1(new_n372), .B2(KEYINPUT31), .ZN(new_n373));
  AOI211_X1 g187(.A(KEYINPUT70), .B(new_n331), .C1(new_n330), .C2(new_n341), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n260), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n368), .A2(new_n260), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT74), .B1(new_n366), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n317), .B1(new_n327), .B2(new_n297), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n333), .A2(KEYINPUT73), .A3(new_n386), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n321), .A2(KEYINPUT73), .A3(new_n332), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n344), .B1(new_n389), .B2(new_n343), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n253), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n330), .A2(new_n348), .A3(new_n333), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n347), .A2(new_n339), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G472), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n385), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n259), .B1(new_n380), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G221), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(new_n253), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT3), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT3), .A2(G107), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(G104), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(KEYINPUT81), .A2(G104), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT81), .A2(G104), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(G104), .B2(G107), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n354), .A2(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n265), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n272), .B2(new_n273), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n326), .B2(new_n268), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n422), .A2(new_n423), .B1(new_n424), .B2(new_n418), .ZN(new_n425));
  INV_X1    g239(.A(new_n411), .ZN(new_n426));
  NOR2_X1   g240(.A1(KEYINPUT81), .A2(G104), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n426), .A2(new_n427), .A3(new_n405), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT3), .A2(G107), .ZN(new_n429));
  INV_X1    g243(.A(G104), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n410), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n414), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(G101), .C1(new_n428), .C2(new_n431), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n320), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT82), .ZN(new_n437));
  INV_X1    g251(.A(new_n319), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n433), .A2(new_n439), .A3(new_n320), .A4(new_n435), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n425), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G140), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n237), .A2(G227), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n324), .A2(new_n325), .B1(new_n419), .B2(new_n265), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n414), .A2(new_n417), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n423), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n418), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n440), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n438), .B1(new_n450), .B2(new_n437), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n444), .B(KEYINPUT80), .Z(new_n453));
  NOR2_X1   g267(.A1(new_n418), .A2(new_n274), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n446), .A2(new_n447), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n319), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n356), .A2(new_n447), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n438), .B1(new_n422), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT12), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n453), .B1(new_n462), .B2(new_n441), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n452), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n460), .A2(KEYINPUT12), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n457), .B(new_n438), .C1(new_n422), .C2(new_n459), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n441), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n453), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  INV_X1    g284(.A(new_n437), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n440), .A2(new_n448), .A3(new_n449), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n319), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n441), .A3(new_n444), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n464), .A2(G469), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n465), .A2(new_n466), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n445), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n444), .B1(new_n473), .B2(new_n441), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n253), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n477), .A2(new_n253), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n403), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n433), .A2(new_n317), .A3(new_n435), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n313), .A2(new_n314), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT5), .A3(new_n299), .ZN(new_n490));
  OAI21_X1  g304(.A(G113), .B1(new_n299), .B2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n418), .A2(new_n316), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G122), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n494), .A3(new_n496), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n326), .A2(new_n209), .A3(new_n268), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n294), .A2(G125), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G224), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(G953), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n495), .A2(new_n510), .A3(new_n497), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n500), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n496), .B(KEYINPUT8), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n491), .B1(new_n315), .B2(KEYINPUT5), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n489), .A2(new_n299), .A3(new_n309), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n447), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n493), .A2(new_n316), .B1(new_n414), .B2(new_n417), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n503), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n499), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n506), .B2(new_n508), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n513), .B(new_n253), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n526), .A2(new_n527), .B1(KEYINPUT7), .B2(new_n505), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n499), .A3(new_n519), .A4(new_n521), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n513), .B1(new_n529), .B2(new_n253), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n487), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n253), .B1(new_n522), .B2(new_n523), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(new_n486), .A3(new_n512), .A4(new_n524), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G237), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n237), .A3(G214), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n263), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n335), .A2(G143), .A3(G214), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n280), .A3(new_n539), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n280), .B1(new_n538), .B2(new_n539), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n544), .A2(new_n215), .A3(new_n216), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n539), .ZN(new_n548));
  AOI21_X1  g362(.A(G143), .B1(new_n335), .B2(G214), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(KEYINPUT18), .A2(G131), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n208), .A2(new_n210), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G146), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n550), .A2(new_n552), .B1(new_n233), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n551), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT86), .B1(new_n540), .B2(new_n551), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n430), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n547), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n547), .B2(new_n559), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT90), .B(new_n253), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n547), .A2(new_n559), .ZN(new_n567));
  INV_X1    g381(.A(new_n561), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n562), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT90), .B1(new_n570), .B2(new_n253), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n233), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n232), .A2(new_n214), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n575), .A2(new_n576), .B1(new_n540), .B2(new_n551), .ZN(new_n577));
  INV_X1    g391(.A(new_n558), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(new_n556), .ZN(new_n579));
  INV_X1    g393(.A(new_n543), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n545), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n208), .A2(new_n210), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n214), .C1(new_n584), .C2(new_n232), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n230), .A2(new_n231), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n581), .B1(new_n586), .B2(KEYINPUT88), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT88), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n230), .A2(new_n588), .A3(new_n585), .A4(new_n231), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n579), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n561), .B1(new_n590), .B2(KEYINPUT89), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(KEYINPUT88), .ZN(new_n592));
  INV_X1    g406(.A(new_n581), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n559), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT89), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n563), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(G475), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n574), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n559), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n568), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n590), .A2(KEYINPUT89), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n562), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n599), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n572), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G478), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n610));
  AND2_X1   g424(.A1(KEYINPUT91), .A2(G122), .ZN(new_n611));
  NOR2_X1   g425(.A1(KEYINPUT91), .A2(G122), .ZN(new_n612));
  OAI21_X1  g426(.A(G116), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n301), .A2(G122), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n409), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n263), .A2(G128), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G134), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n276), .A3(new_n617), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  INV_X1    g436(.A(new_n612), .ZN(new_n623));
  NAND2_X1  g437(.A1(KEYINPUT91), .A2(G122), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n301), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(G122), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT14), .B1(new_n626), .B2(G116), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT14), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n301), .A3(G122), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n622), .B(G107), .C1(new_n625), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n613), .A2(new_n627), .A3(new_n629), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n622), .B1(new_n633), .B2(G107), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n615), .B(new_n621), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n614), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G107), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n615), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT13), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n616), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n618), .A3(G134), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n616), .B(new_n617), .C1(new_n639), .C2(new_n276), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n400), .A2(new_n256), .A3(G953), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n635), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n635), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n253), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n635), .A2(new_n643), .ZN(new_n650));
  INV_X1    g464(.A(new_n644), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n635), .A2(new_n643), .A3(new_n644), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(KEYINPUT94), .A3(new_n253), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n610), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n648), .B(G902), .C1(new_n652), .C2(new_n653), .ZN(new_n657));
  INV_X1    g471(.A(new_n610), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(G234), .A2(G237), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(G952), .A3(new_n237), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(G902), .A3(G953), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT21), .B(G898), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n656), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(G214), .B1(G237), .B2(G902), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n535), .A2(new_n608), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT95), .B1(new_n485), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n535), .A2(new_n667), .A3(new_n668), .ZN(new_n671));
  INV_X1    g485(.A(new_n444), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n438), .A2(new_n425), .A3(new_n437), .A4(new_n440), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n451), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n462), .A2(new_n441), .A3(new_n444), .ZN(new_n675));
  AOI21_X1  g489(.A(G902), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n482), .B1(new_n676), .B2(new_n477), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n464), .A2(G469), .A3(new_n475), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n402), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT95), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n671), .A2(new_n679), .A3(new_n680), .A4(new_n608), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n670), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n398), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n413), .ZN(G3));
  AND2_X1   g498(.A1(new_n679), .A2(new_n259), .ZN(new_n685));
  INV_X1    g499(.A(new_n608), .ZN(new_n686));
  INV_X1    g500(.A(G478), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n647), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT96), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n654), .B(KEYINPUT33), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(G478), .A3(new_n253), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n668), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n531), .B2(new_n534), .ZN(new_n696));
  INV_X1    g510(.A(new_n666), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n366), .B2(G902), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n377), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n685), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT97), .Z(new_n704));
  XOR2_X1   g518(.A(KEYINPUT34), .B(G104), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G6));
  INV_X1    g520(.A(KEYINPUT98), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n598), .A2(new_n600), .A3(new_n574), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n573), .B1(new_n605), .B2(new_n599), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n605), .A2(new_n599), .A3(new_n573), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n601), .A2(new_n711), .A3(KEYINPUT98), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT94), .B1(new_n654), .B2(new_n253), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n658), .B1(new_n713), .B2(new_n657), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n655), .A2(new_n610), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n572), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n698), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n685), .A2(new_n702), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT35), .B(G107), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G9));
  NOR2_X1   g535(.A1(new_n249), .A2(new_n250), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n246), .A2(KEYINPUT36), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n701), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n670), .A2(new_n681), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT37), .B(G110), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G12));
  AOI21_X1  g543(.A(KEYINPUT25), .B1(new_n252), .B2(new_n253), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n187), .B(G902), .C1(new_n251), .C2(new_n240), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n257), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n258), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n679), .B(new_n734), .C1(new_n380), .C2(new_n397), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n601), .A2(KEYINPUT98), .A3(new_n711), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT98), .B1(new_n601), .B2(new_n711), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n661), .B(KEYINPUT99), .Z(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(G900), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n664), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n739), .A2(KEYINPUT100), .A3(new_n716), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n710), .A2(new_n716), .A3(new_n712), .A4(new_n744), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n696), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT101), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT101), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n748), .A3(new_n751), .A4(new_n696), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n736), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G128), .ZN(G30));
  XOR2_X1   g568(.A(new_n743), .B(KEYINPUT39), .Z(new_n755));
  NAND2_X1  g569(.A1(new_n679), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT40), .Z(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n535), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n656), .A2(new_n659), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n686), .A2(new_n761), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n759), .A2(new_n734), .A3(new_n762), .A4(new_n695), .ZN(new_n763));
  INV_X1    g577(.A(new_n389), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n253), .B1(new_n764), .B2(new_n339), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n348), .B1(new_n330), .B2(new_n333), .ZN(new_n766));
  OAI21_X1  g580(.A(G472), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n383), .A2(new_n385), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n757), .B(new_n763), .C1(new_n380), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT103), .B(G143), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G45));
  NOR3_X1   g585(.A1(new_n366), .A2(KEYINPUT74), .A3(new_n382), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n384), .B1(new_n375), .B2(new_n381), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n370), .A3(new_n379), .A4(new_n396), .ZN(new_n775));
  INV_X1    g589(.A(new_n696), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n694), .A2(new_n776), .A3(new_n743), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n679), .A3(new_n734), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G146), .ZN(G48));
  NOR2_X1   g593(.A1(new_n479), .A2(new_n480), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n780), .B2(G902), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n403), .A3(new_n481), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n775), .A2(new_n259), .A3(new_n699), .A4(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT41), .B(G113), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT104), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n784), .B(new_n786), .ZN(G15));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n259), .A3(new_n718), .A4(new_n783), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G116), .ZN(G18));
  NOR2_X1   g603(.A1(new_n669), .A2(new_n782), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n775), .A2(new_n734), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G119), .ZN(G21));
  NAND2_X1  g606(.A1(new_n390), .A2(new_n348), .ZN(new_n793));
  INV_X1    g607(.A(new_n363), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT105), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n342), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n793), .B2(new_n794), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n376), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n700), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n762), .A2(new_n666), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n776), .A2(new_n782), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n259), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G122), .ZN(G24));
  AND3_X1   g618(.A1(new_n734), .A2(new_n799), .A3(new_n700), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n694), .A2(new_n743), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n802), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT106), .B(G125), .Z(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G27));
  OAI211_X1 g623(.A(new_n369), .B(new_n396), .C1(new_n366), .C2(new_n382), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n259), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n469), .A2(G469), .A3(new_n474), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n481), .A2(new_n483), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n403), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n531), .A2(new_n668), .A3(new_n534), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT107), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n531), .A2(new_n668), .A3(new_n534), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT107), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n819), .A3(new_n403), .A4(new_n814), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n812), .A2(KEYINPUT42), .A3(new_n806), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n775), .A2(new_n259), .A3(new_n806), .A4(new_n821), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT108), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT42), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n823), .B2(KEYINPUT108), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G131), .ZN(G33));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n748), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n775), .A3(new_n259), .A4(new_n821), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n746), .B(KEYINPUT100), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT109), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n821), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n398), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  INV_X1    g651(.A(new_n745), .ZN(new_n838));
  INV_X1    g652(.A(new_n748), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(KEYINPUT110), .A3(new_n840), .A4(new_n830), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G134), .ZN(G36));
  AOI21_X1  g657(.A(KEYINPUT45), .B1(new_n464), .B2(new_n475), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n469), .A2(KEYINPUT45), .A3(new_n474), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(G469), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n483), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT46), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n847), .A2(new_n848), .B1(new_n477), .B2(new_n676), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n402), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n755), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n693), .A2(new_n608), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT43), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT43), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n693), .A2(new_n855), .A3(new_n608), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n701), .A3(new_n734), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT44), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n816), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n852), .B(new_n859), .C1(new_n858), .C2(new_n857), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(G137), .ZN(G39));
  INV_X1    g675(.A(KEYINPUT111), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT47), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n851), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n806), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n775), .A2(new_n865), .A3(new_n259), .A4(new_n816), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n862), .A2(KEYINPUT47), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n851), .B1(new_n867), .B2(new_n863), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(G140), .ZN(G42));
  NAND2_X1  g684(.A1(new_n781), .A2(new_n481), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n402), .B(new_n695), .C1(new_n871), .C2(KEYINPUT49), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(KEYINPUT49), .B2(new_n871), .ZN(new_n873));
  INV_X1    g687(.A(new_n759), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n853), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n380), .A2(new_n768), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n259), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n854), .A2(new_n741), .A3(new_n856), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n879), .A2(new_n259), .A3(new_n800), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n695), .A3(new_n759), .A4(new_n783), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT50), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n783), .A2(new_n818), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT115), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n259), .A2(new_n884), .A3(new_n662), .A4(new_n876), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n608), .A2(new_n690), .A3(new_n692), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n884), .A2(new_n879), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n885), .A2(new_n887), .B1(new_n805), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n871), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n402), .B1(new_n890), .B2(KEYINPUT114), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(KEYINPUT114), .B2(new_n890), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n864), .B2(new_n868), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n880), .A2(new_n818), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n882), .B(new_n889), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n752), .A2(new_n775), .A3(new_n679), .A4(new_n734), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n751), .B1(new_n832), .B2(new_n696), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n734), .A2(new_n743), .A3(new_n815), .ZN(new_n905));
  AND4_X1   g719(.A1(new_n686), .A2(new_n668), .A3(new_n535), .A4(new_n761), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n380), .C2(new_n768), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n778), .A2(new_n807), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n778), .A2(new_n807), .A3(new_n907), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(new_n910), .B2(new_n753), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n784), .A2(new_n788), .A3(new_n791), .A4(new_n803), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n694), .B1(new_n686), .B2(new_n760), .ZN(new_n914));
  INV_X1    g728(.A(new_n698), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n685), .A2(new_n914), .A3(new_n915), .A4(new_n702), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n727), .B(new_n916), .C1(new_n398), .C2(new_n682), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n821), .A2(new_n805), .A3(new_n806), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n761), .A2(new_n572), .A3(new_n743), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n739), .A3(new_n818), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n735), .B2(new_n920), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n913), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n827), .A3(new_n842), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n900), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n822), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n775), .A2(new_n259), .A3(new_n806), .A4(new_n821), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT108), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT42), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n823), .A2(KEYINPUT108), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n917), .A2(new_n921), .ZN(new_n931));
  AND4_X1   g745(.A1(new_n784), .A2(new_n788), .A3(new_n791), .A4(new_n803), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n904), .B1(new_n903), .B2(new_n908), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n910), .A2(KEYINPUT52), .A3(new_n753), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n934), .A2(KEYINPUT53), .A3(new_n842), .A4(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n924), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n912), .B2(new_n923), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n943));
  OR3_X1    g757(.A1(new_n912), .A2(new_n923), .A3(new_n900), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT112), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(new_n941), .C1(new_n912), .C2(new_n923), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n947), .B2(KEYINPUT54), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n885), .A2(new_n686), .A3(new_n693), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n237), .A2(G952), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n880), .B2(new_n802), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT48), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n888), .A2(new_n952), .A3(new_n812), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n888), .B2(new_n812), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n949), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n895), .B2(new_n896), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n899), .A2(new_n948), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n877), .B1(new_n957), .B2(new_n958), .ZN(G75));
  NOR2_X1   g773(.A1(new_n237), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n253), .B1(new_n924), .B2(new_n938), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(G210), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT56), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n500), .A2(new_n511), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(new_n509), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n968), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT117), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n965), .A2(KEYINPUT117), .A3(new_n968), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G51));
  NAND2_X1  g788(.A1(new_n924), .A2(new_n938), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT54), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n924), .A2(new_n938), .A3(new_n939), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n482), .B(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n780), .B(KEYINPUT118), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n844), .A2(new_n846), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n962), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n960), .B1(new_n982), .B2(new_n984), .ZN(G54));
  NAND3_X1  g799(.A1(new_n962), .A2(KEYINPUT58), .A3(G475), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n960), .B1(new_n986), .B2(new_n598), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n598), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT119), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT119), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n987), .B(new_n990), .C1(new_n598), .C2(new_n986), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G60));
  INV_X1    g806(.A(KEYINPUT122), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n691), .B(KEYINPUT120), .ZN(new_n994));
  XNOR2_X1  g808(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n687), .A2(new_n253), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n993), .B1(new_n978), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n939), .B1(new_n924), .B2(new_n938), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n993), .B(new_n998), .C1(new_n940), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n961), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n948), .B2(new_n997), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT123), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT123), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1006), .B(new_n994), .C1(new_n948), .C2(new_n997), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n1005), .B2(new_n1007), .ZN(G63));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT60), .Z(new_n1010));
  NAND3_X1  g824(.A1(new_n975), .A2(new_n724), .A3(new_n1010), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n975), .A2(new_n1010), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n252), .B(KEYINPUT124), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n961), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g829(.A(G953), .B1(new_n665), .B2(new_n504), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n913), .A2(new_n917), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n966), .B1(G898), .B2(new_n237), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT125), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1018), .B(new_n1020), .ZN(G69));
  NOR2_X1   g835(.A1(new_n584), .A2(new_n232), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n232), .B2(new_n582), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n360), .B(new_n1023), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n753), .A2(new_n778), .A3(new_n807), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n769), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n756), .A2(new_n816), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1028), .A2(new_n775), .A3(new_n259), .A4(new_n914), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n860), .A2(new_n869), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1024), .B1(new_n1032), .B2(new_n237), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1024), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n742), .A2(new_n237), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1025), .A2(new_n842), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n852), .A2(new_n812), .A3(new_n906), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n860), .A2(new_n869), .A3(new_n1037), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n1036), .A2(new_n1038), .A3(new_n930), .ZN(new_n1039));
  AOI211_X1 g853(.A(new_n1034), .B(new_n1035), .C1(new_n1039), .C2(new_n237), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n237), .B1(G227), .B2(G900), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1042), .A2(KEYINPUT126), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1033), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1042), .A2(KEYINPUT126), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1044), .B(new_n1045), .Z(G72));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  INV_X1    g862(.A(new_n1017), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1048), .B1(new_n1032), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n960), .B1(new_n1050), .B2(new_n766), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1039), .A2(new_n1017), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT127), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1052), .A2(new_n1053), .A3(new_n1048), .ZN(new_n1054));
  INV_X1    g868(.A(new_n393), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1052), .B2(new_n1048), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1051), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1048), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1055), .A2(new_n766), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1058), .B1(new_n947), .B2(new_n1060), .ZN(G57));
endmodule


