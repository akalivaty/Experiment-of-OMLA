//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G250), .B(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G264), .B(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n229), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G45), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n243), .A2(G1), .ZN(new_n244));
  INV_X1    g0044(.A(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT5), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G270), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT78), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n247), .B2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n245), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n256));
  AND4_X1   g0056(.A1(new_n255), .A2(new_n256), .A3(new_n244), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(G274), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT79), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n255), .A2(new_n256), .A3(new_n244), .A4(new_n248), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT79), .B1(new_n262), .B2(new_n258), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n253), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n251), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(G257), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G303), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n273), .A2(G264), .A3(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n265), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n264), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n284), .A3(KEYINPUT68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  INV_X1    g0086(.A(G20), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n282), .A2(new_n287), .A3(G1), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n285), .A2(new_n289), .A3(G116), .A4(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G116), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(G20), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G283), .ZN(new_n295));
  INV_X1    g0095(.A(G97), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n287), .C1(G33), .C2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n280), .C1(new_n287), .C2(G116), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT20), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n292), .B(new_n294), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n277), .A2(new_n302), .A3(KEYINPUT21), .A4(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT82), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n264), .B2(new_n276), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT82), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT21), .A4(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n277), .B2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n277), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT21), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n264), .A2(G179), .A3(new_n276), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n313), .A2(new_n314), .B1(new_n316), .B2(new_n302), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n309), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT8), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(G58), .ZN(new_n320));
  INV_X1    g0120(.A(G58), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(KEYINPUT8), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT67), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(KEYINPUT8), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(G58), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(new_n287), .A3(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G20), .A2(G33), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n281), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n288), .A2(new_n202), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n290), .A2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(new_n279), .A3(new_n278), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n202), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n273), .A2(G222), .A3(new_n270), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n273), .A2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G223), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n339), .B1(new_n340), .B2(new_n273), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n265), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT66), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n290), .C1(G41), .C2(G45), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n251), .A3(G274), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n245), .A2(new_n243), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n290), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n290), .A2(new_n349), .B1(new_n210), .B2(new_n250), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(G226), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n344), .A2(new_n353), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n305), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n338), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n332), .B2(new_n336), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n344), .A2(G190), .A3(new_n353), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  INV_X1    g0163(.A(new_n336), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n329), .A2(new_n331), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT9), .B(new_n364), .C1(new_n365), .C2(new_n281), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(G200), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n362), .A2(new_n363), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n366), .A2(new_n361), .A3(new_n360), .A4(new_n367), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n358), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n285), .A2(new_n289), .A3(G77), .A4(new_n334), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT8), .B(G58), .ZN(new_n373));
  INV_X1    g0173(.A(new_n330), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n287), .B2(new_n340), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n287), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n280), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n372), .B(new_n379), .C1(G77), .C2(new_n284), .ZN(new_n380));
  INV_X1    g0180(.A(G107), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n341), .A2(new_n216), .B1(new_n381), .B2(new_n273), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n267), .A2(new_n269), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n383), .A2(new_n231), .A3(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n265), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n351), .B1(G244), .B2(new_n352), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n388), .B2(G169), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(G179), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT69), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n388), .A2(new_n393), .B1(new_n394), .B2(new_n380), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n380), .A2(new_n394), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n311), .B2(new_n387), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n371), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n383), .B2(new_n287), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n402), .B(G20), .C1(new_n267), .C2(new_n269), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(G58), .C2(G68), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(G20), .B1(G159), .B2(new_n330), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n273), .B2(G20), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n268), .A2(G33), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT7), .B(new_n287), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n215), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n330), .A2(G159), .ZN(new_n417));
  INV_X1    g0217(.A(new_n407), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n418), .A2(new_n405), .A3(new_n201), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n287), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n411), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n410), .A2(new_n421), .A3(new_n280), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n284), .B1(new_n323), .B2(new_n327), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n373), .A2(new_n324), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT67), .B1(new_n320), .B2(new_n322), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n335), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT74), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n423), .B2(new_n426), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n347), .A2(new_n251), .A3(G274), .ZN(new_n433));
  INV_X1    g0233(.A(new_n350), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n433), .A2(new_n434), .B1(G232), .B2(new_n352), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n267), .A2(new_n269), .A3(G226), .A4(G1698), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n267), .A2(new_n269), .A3(G223), .A4(new_n270), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n265), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(new_n345), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n290), .B1(G41), .B2(G45), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n251), .A2(G232), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n348), .B2(new_n350), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n265), .B2(new_n439), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n441), .B1(new_n445), .B2(G169), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n431), .A2(new_n432), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n432), .B1(new_n431), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT75), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n424), .A2(new_n425), .A3(new_n335), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n288), .B1(new_n424), .B2(new_n425), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT74), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n423), .A2(new_n427), .A3(new_n426), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n404), .A2(new_n409), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n281), .B1(new_n456), .B2(new_n411), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n457), .B2(new_n410), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT18), .B1(new_n458), .B2(new_n446), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n446), .B1(new_n422), .B2(new_n430), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n432), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n435), .A2(new_n440), .A3(new_n311), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n445), .B2(G200), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n422), .A2(new_n465), .A3(new_n430), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n422), .A2(new_n465), .A3(new_n430), .A4(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n450), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n433), .A2(new_n434), .B1(G238), .B2(new_n352), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n267), .A2(new_n269), .A3(G232), .A4(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n267), .A2(new_n269), .A3(G226), .A4(new_n270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G97), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n265), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT13), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n473), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n473), .B2(new_n478), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT14), .B1(new_n482), .B2(new_n305), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT14), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(G169), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT72), .B1(new_n482), .B2(G179), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT72), .ZN(new_n487));
  NOR4_X1   g0287(.A1(new_n480), .A2(new_n481), .A3(new_n487), .A4(new_n345), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n284), .B2(G68), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n284), .A2(new_n490), .A3(G68), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT12), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n490), .B(KEYINPUT12), .C1(new_n284), .C2(G68), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n330), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n340), .B2(new_n377), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n280), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT11), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n285), .A2(new_n289), .A3(G68), .A4(new_n334), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n503));
  AND4_X1   g0303(.A1(new_n496), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n489), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n481), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n473), .A2(new_n478), .A3(new_n479), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(G190), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G200), .B1(new_n480), .B2(new_n481), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n504), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n509), .A2(new_n510), .A3(new_n504), .A4(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n400), .A2(new_n472), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n267), .A2(new_n269), .A3(G257), .A4(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n267), .A2(new_n269), .A3(G250), .A4(new_n270), .ZN(new_n519));
  INV_X1    g0319(.A(G294), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n519), .C1(new_n266), .C2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n261), .A2(new_n263), .B1(new_n521), .B2(new_n265), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n249), .A2(G264), .A3(new_n251), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(KEYINPUT86), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT86), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n249), .A2(new_n526), .A3(G264), .A4(new_n251), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n524), .A2(new_n305), .B1(new_n345), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT23), .B1(new_n287), .B2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n381), .A3(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n287), .A2(G33), .A3(G116), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT83), .A2(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n273), .A2(new_n287), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n273), .A2(KEYINPUT22), .A3(new_n287), .A4(new_n538), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n280), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n288), .A2(new_n280), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n291), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT25), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n284), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n381), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n550), .A2(G107), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT85), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n539), .A2(new_n540), .ZN(new_n557));
  INV_X1    g0357(.A(new_n537), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n543), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n542), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n281), .B1(new_n561), .B2(new_n544), .ZN(new_n562));
  INV_X1    g0362(.A(new_n554), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n530), .A2(new_n555), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n267), .A2(new_n269), .A3(G238), .A4(new_n270), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n267), .A2(new_n269), .A3(G244), .A4(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n265), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n218), .B1(new_n243), .B2(G1), .ZN(new_n571));
  INV_X1    g0371(.A(G274), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n290), .A2(new_n572), .A3(G45), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n251), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n305), .ZN(new_n576));
  NAND3_X1  g0376(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(new_n287), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G87), .A2(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n381), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(KEYINPUT80), .A3(new_n381), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n267), .A2(new_n269), .A3(new_n287), .A4(G68), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n377), .B2(new_n296), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n280), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n376), .A2(new_n288), .ZN(new_n590));
  INV_X1    g0390(.A(new_n376), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n548), .A2(new_n291), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n574), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n569), .B2(new_n265), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n345), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n576), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n548), .A2(G87), .A3(new_n291), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n589), .A2(new_n599), .A3(new_n590), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n595), .A2(new_n393), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n311), .B(new_n594), .C1(new_n569), .C2(new_n265), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT81), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n602), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n589), .A2(new_n590), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n575), .A2(G200), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n599), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT81), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n597), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n522), .A2(new_n311), .A3(new_n523), .ZN(new_n612));
  AOI21_X1  g0412(.A(G200), .B1(new_n522), .B2(new_n528), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n547), .B(new_n554), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n288), .A2(new_n296), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(KEYINPUT76), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n549), .C2(new_n296), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n330), .A2(G77), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT6), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n620), .A2(new_n296), .A3(G107), .ZN(new_n621));
  XNOR2_X1  g0421(.A(G97), .B(G107), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n623), .B2(new_n287), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n381), .B1(new_n412), .B2(new_n415), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n618), .B1(new_n626), .B2(new_n280), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n267), .A2(new_n269), .A3(G244), .A4(new_n270), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT77), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT4), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n273), .A2(G244), .A3(new_n270), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n631), .A2(new_n295), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n265), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n249), .A2(G257), .A3(new_n251), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n261), .B2(new_n263), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n636), .A2(new_n639), .A3(new_n311), .ZN(new_n640));
  AOI21_X1  g0440(.A(G200), .B1(new_n636), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n627), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n636), .A2(new_n639), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n305), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n280), .B1(new_n624), .B2(new_n625), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n550), .A2(G97), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n616), .A4(new_n617), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n636), .A2(new_n639), .A3(new_n345), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n614), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n318), .A2(new_n517), .A3(new_n565), .A4(new_n651), .ZN(G372));
  AND2_X1   g0452(.A1(new_n489), .A2(new_n505), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n391), .B1(new_n513), .B2(new_n514), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT89), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n515), .A2(new_n392), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n506), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n658), .A3(new_n471), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n459), .A2(new_n461), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n368), .A2(new_n370), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n358), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n611), .B2(new_n649), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT87), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n606), .A2(new_n607), .A3(new_n666), .A4(new_n599), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT87), .B1(new_n600), .B2(new_n601), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n605), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n597), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  INV_X1    g0472(.A(new_n649), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n597), .B(KEYINPUT88), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n665), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n530), .B1(new_n562), .B2(new_n563), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n309), .A3(new_n317), .ZN(new_n678));
  INV_X1    g0478(.A(new_n650), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n671), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n517), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n664), .A2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n283), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .A3(G20), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT27), .B1(new_n685), .B2(G20), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n302), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n318), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n309), .A2(new_n317), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n302), .A3(new_n690), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n684), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n565), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n690), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n555), .A2(new_n564), .A3(new_n690), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n565), .A2(new_n698), .A3(new_n614), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n690), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n699), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n677), .A2(new_n690), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n701), .A2(new_n706), .ZN(G399));
  NAND3_X1  g0507(.A1(new_n582), .A2(new_n293), .A3(new_n583), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n207), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n213), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n565), .A2(new_n309), .A3(new_n317), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(new_n679), .A3(new_n671), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT26), .B1(new_n670), .B2(new_n649), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n604), .A2(new_n673), .A3(new_n672), .A4(new_n610), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n675), .A3(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n702), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n690), .B1(new_n676), .B2(new_n680), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n651), .A2(new_n318), .A3(new_n565), .A4(new_n702), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n636), .A2(new_n639), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n525), .A2(new_n527), .B1(new_n521), .B2(new_n265), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(new_n595), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n316), .A2(new_n725), .A3(new_n727), .A4(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n636), .A2(new_n726), .A3(new_n639), .A4(new_n595), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n315), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n595), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n529), .A2(new_n643), .A3(new_n277), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n734), .B2(new_n690), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n723), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n715), .B1(new_n741), .B2(G1), .ZN(G364));
  NOR2_X1   g0542(.A1(new_n282), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n290), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n711), .A2(new_n745), .A3(KEYINPUT90), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT90), .B1(new_n711), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n695), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n692), .A2(new_n694), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(G330), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n279), .B1(G20), .B2(new_n305), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n287), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n393), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n273), .B1(new_n757), .B2(new_n381), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n287), .A2(new_n311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n345), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n755), .A2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G58), .A2(new_n762), .B1(new_n764), .B2(G77), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(KEYINPUT92), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT32), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n758), .B(new_n767), .C1(new_n768), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n287), .B1(new_n769), .B2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n296), .ZN(new_n775));
  NAND3_X1  g0575(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n311), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n772), .A2(new_n768), .B1(new_n202), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n776), .A2(G190), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n775), .B(new_n779), .C1(G68), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(KEYINPUT92), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n759), .A2(new_n756), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n773), .A2(new_n781), .A3(new_n782), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(G303), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n383), .B1(new_n757), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n780), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n774), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G294), .B1(G326), .B2(new_n777), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n761), .A2(new_n797), .B1(new_n763), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n770), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G329), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n790), .A2(new_n794), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n754), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G13), .A2(G33), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G20), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n753), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n273), .A2(new_n207), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT91), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(G116), .B2(new_n207), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n710), .A2(new_n273), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G45), .B2(new_n213), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n241), .B2(G45), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n748), .B(new_n803), .C1(new_n807), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n806), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n751), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n752), .A2(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n391), .A2(new_n690), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n380), .A2(new_n690), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n395), .C2(new_n397), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n391), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n722), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n749), .B1(new_n826), .B2(new_n739), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n739), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n757), .A2(new_n217), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G116), .B2(new_n764), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n830), .B1(new_n520), .B2(new_n761), .C1(new_n786), .C2(new_n381), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n383), .B1(new_n770), .B2(new_n798), .ZN(new_n832));
  INV_X1    g0632(.A(new_n780), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n833), .A2(new_n791), .B1(new_n778), .B2(new_n272), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n831), .A2(new_n775), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT94), .Z(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n762), .B1(new_n764), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n833), .B2(new_n838), .C1(new_n839), .C2(new_n778), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n787), .A2(G50), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n774), .A2(new_n321), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n273), .B1(new_n757), .B2(new_n215), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G132), .C2(new_n800), .ZN(new_n847));
  AND4_X1   g0647(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n753), .B1(new_n836), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n753), .A2(new_n804), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n748), .B1(new_n340), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n825), .C2(new_n805), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n828), .A2(new_n852), .ZN(G384));
  NAND2_X1  g0653(.A1(new_n622), .A2(new_n620), .ZN(new_n854));
  INV_X1    g0654(.A(new_n621), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(new_n293), .A4(new_n212), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  OR4_X1    g0660(.A1(new_n340), .A2(new_n418), .A3(new_n213), .A4(new_n405), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n202), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n290), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n431), .A2(new_n447), .ZN(new_n865));
  INV_X1    g0665(.A(new_n688), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n431), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n867), .A3(new_n466), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT96), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n865), .A2(new_n867), .A3(new_n871), .A4(new_n466), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n472), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n422), .A2(new_n465), .A3(new_n430), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n460), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n871), .B1(new_n881), .B2(new_n867), .ZN(new_n882));
  AND4_X1   g0682(.A1(new_n871), .A2(new_n865), .A3(new_n867), .A4(new_n466), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT96), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND4_X1   g0684(.A1(KEYINPUT38), .A2(new_n877), .A3(new_n879), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .A4(new_n884), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n867), .B1(new_n661), .B2(new_n471), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n882), .A2(new_n883), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(KEYINPUT98), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n506), .A2(new_n690), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n884), .A2(new_n879), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n470), .B1(new_n660), .B2(KEYINPUT75), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n867), .B1(new_n897), .B2(new_n463), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n887), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT98), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n894), .A2(new_n895), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n505), .A2(new_n690), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n506), .A2(new_n515), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n506), .B2(new_n515), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n665), .A2(new_n674), .A3(new_n675), .ZN(new_n909));
  INV_X1    g0709(.A(new_n680), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n702), .B(new_n825), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n820), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n900), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n660), .A2(new_n688), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT97), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT97), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n903), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n517), .B(new_n721), .C1(new_n722), .C2(KEYINPUT29), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n664), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT99), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n724), .A2(new_n737), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n825), .B1(new_n905), .B2(new_n906), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n724), .B2(new_n737), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n900), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n887), .B2(new_n892), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n929), .A2(new_n930), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n738), .A2(KEYINPUT99), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n724), .A2(new_n737), .A3(new_n924), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n517), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(G330), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n923), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n290), .B2(new_n743), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n923), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n864), .B1(new_n941), .B2(new_n942), .ZN(G367));
  INV_X1    g0743(.A(KEYINPUT103), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n649), .B(new_n642), .C1(new_n627), .C2(new_n702), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT100), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT100), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n673), .A2(new_n690), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n704), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n950), .A2(KEYINPUT42), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT42), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n946), .A2(new_n947), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n673), .B1(new_n954), .B2(new_n696), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n952), .B(new_n953), .C1(new_n690), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n600), .A2(new_n690), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n671), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n675), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n956), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n962), .B1(new_n956), .B2(new_n963), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n965), .A2(new_n966), .B1(new_n701), .B2(new_n950), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n701), .A2(new_n950), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n711), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n706), .A2(new_n949), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n706), .A2(new_n949), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n701), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n701), .B1(new_n975), .B2(new_n977), .ZN(new_n980));
  INV_X1    g0780(.A(new_n703), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n951), .B1(new_n700), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n695), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n741), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n973), .B1(new_n985), .B2(new_n740), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n971), .B1(new_n986), .B2(new_n744), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n807), .B1(new_n207), .B2(new_n376), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n228), .B2(new_n812), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n786), .A2(new_n321), .B1(new_n839), .B2(new_n770), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT102), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n383), .B1(new_n762), .B2(G150), .ZN(new_n992));
  INV_X1    g0792(.A(new_n757), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G50), .A2(new_n764), .B1(new_n993), .B2(G77), .ZN(new_n994));
  INV_X1    g0794(.A(G143), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n833), .A2(new_n771), .B1(new_n778), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G68), .B2(new_n795), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n991), .A2(new_n992), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n990), .A2(KEYINPUT102), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n786), .A2(new_n293), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT46), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(KEYINPUT101), .B(G317), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n383), .B1(new_n770), .B2(new_n1002), .C1(new_n778), .C2(new_n798), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n833), .A2(new_n520), .B1(new_n774), .B2(new_n381), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G97), .A2(new_n993), .B1(new_n764), .B2(G283), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n272), .C2(new_n761), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n748), .B(new_n989), .C1(new_n1009), .C2(new_n753), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n958), .A2(new_n959), .A3(new_n806), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n944), .B1(new_n987), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n980), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n984), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n978), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n741), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n745), .B1(new_n1018), .B2(new_n973), .ZN(new_n1019));
  OAI211_X1 g0819(.A(KEYINPUT103), .B(new_n1012), .C1(new_n1019), .C2(new_n971), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1014), .A2(new_n1020), .ZN(G387));
  NAND2_X1  g0821(.A1(new_n983), .A2(new_n745), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n812), .B1(new_n234), .B2(new_n243), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n709), .B2(new_n809), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n373), .A2(new_n1025), .A3(G50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n373), .B2(G50), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n709), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1024), .A2(new_n1029), .B1(new_n381), .B2(new_n710), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n807), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n749), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT105), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n787), .A2(G77), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n774), .A2(new_n376), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n273), .B1(new_n757), .B2(new_n296), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G159), .C2(new_n777), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n328), .A2(new_n780), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n763), .A2(new_n215), .B1(new_n770), .B2(new_n838), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G50), .B2(new_n762), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n833), .A2(new_n798), .B1(new_n778), .B2(new_n797), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT106), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n761), .A2(new_n1002), .B1(new_n763), .B2(new_n272), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT106), .B2(new_n1042), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n786), .A2(new_n520), .B1(new_n791), .B2(new_n774), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n273), .B1(new_n800), .B2(G326), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n293), .C2(new_n757), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT49), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1041), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1033), .B1(new_n753), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n700), .B2(new_n817), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n984), .A2(new_n711), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n741), .A2(new_n983), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1022), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(G393));
  OAI21_X1  g0860(.A(new_n984), .B1(new_n979), .B2(new_n980), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n1017), .A3(new_n711), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1015), .A2(new_n745), .A3(new_n978), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n807), .B1(new_n296), .B2(new_n207), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n238), .B2(new_n812), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n795), .A2(G77), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n833), .B2(new_n202), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n763), .A2(new_n373), .B1(new_n770), .B2(new_n995), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n383), .A4(new_n829), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n778), .A2(new_n838), .B1(new_n761), .B2(new_n771), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n215), .C2(new_n786), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT107), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n763), .A2(new_n520), .B1(new_n774), .B2(new_n293), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G303), .B2(new_n780), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT108), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n777), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n383), .B1(new_n770), .B2(new_n797), .C1(new_n381), .C2(new_n757), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n787), .B2(G283), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1072), .A2(KEYINPUT107), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1073), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n748), .B(new_n1065), .C1(new_n1083), .C2(new_n753), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n949), .B2(new_n817), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1062), .A2(new_n1063), .A3(new_n1085), .ZN(G390));
  NAND2_X1  g0886(.A1(new_n824), .A2(new_n391), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n912), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n907), .B1(new_n739), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n904), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n516), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n506), .A2(new_n515), .A3(new_n904), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n934), .A2(new_n1093), .A3(G330), .A4(new_n935), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n913), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n934), .A2(G330), .A3(new_n825), .A4(new_n935), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n907), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n702), .B(new_n1087), .C1(new_n717), .C2(new_n720), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n912), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n684), .B(new_n1088), .C1(new_n724), .C2(new_n737), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n908), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n934), .A2(G330), .A3(new_n517), .A4(new_n935), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n664), .A2(new_n921), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n908), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n895), .B1(new_n887), .B2(new_n892), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1101), .A2(new_n908), .ZN(new_n1111));
  AOI211_X1 g0911(.A(KEYINPUT98), .B(new_n888), .C1(new_n899), .C2(new_n887), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n901), .B1(new_n900), .B2(KEYINPUT39), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n893), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n895), .B1(new_n913), .B2(new_n908), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1110), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n894), .A2(new_n902), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1115), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1117), .A2(new_n1118), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1107), .B(new_n1116), .C1(new_n1119), .C2(new_n1094), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1120), .A2(new_n711), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1116), .B1(new_n1119), .B2(new_n1094), .ZN(new_n1122));
  AOI211_X1 g0922(.A(KEYINPUT109), .B(new_n1106), .C1(new_n1096), .C2(new_n1103), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT109), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1106), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1122), .A2(new_n1128), .A3(KEYINPUT110), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT110), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1121), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1122), .A2(new_n744), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n850), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n749), .B1(new_n328), .B2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n778), .A2(new_n791), .B1(new_n763), .B2(new_n296), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G107), .B2(new_n780), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT112), .Z(new_n1137));
  AOI21_X1  g0937(.A(new_n273), .B1(new_n993), .B2(G68), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G116), .A2(new_n762), .B1(new_n800), .B2(G294), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n788), .A2(new_n1066), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OR3_X1    g0940(.A1(new_n786), .A2(KEYINPUT53), .A3(new_n838), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n762), .A2(G132), .B1(new_n764), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n778), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT53), .B1(new_n786), .B2(new_n838), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n795), .A2(G159), .B1(G137), .B2(new_n780), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1141), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n273), .B1(new_n757), .B2(new_n202), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G125), .B2(new_n800), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT111), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1137), .A2(new_n1140), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1134), .B1(new_n1154), .B2(new_n753), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1114), .B2(new_n805), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(G378));
  AOI21_X1  g0958(.A(KEYINPUT97), .B1(new_n914), .B2(new_n915), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1114), .B2(new_n895), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT117), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n663), .A2(new_n357), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT115), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n337), .A2(new_n688), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT55), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n371), .A2(KEYINPUT115), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n371), .A2(KEYINPUT115), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1163), .B(new_n358), .C1(new_n368), .C2(new_n370), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1161), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n932), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n899), .A2(new_n887), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n934), .A2(new_n1093), .A3(new_n935), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n930), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n928), .A2(new_n931), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(G330), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1176), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1160), .A2(new_n1177), .A3(new_n1184), .A4(new_n916), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1176), .B1(new_n932), .B2(G330), .ZN(new_n1186));
  AND4_X1   g0986(.A1(G330), .A2(new_n1180), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n920), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1185), .A2(new_n1188), .A3(KEYINPUT118), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT118), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n711), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n804), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n273), .A2(G41), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G50), .B(new_n1199), .C1(new_n266), .C2(new_n245), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n791), .B2(new_n770), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n757), .A2(new_n321), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1034), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT113), .Z(new_n1205));
  OAI22_X1  g1005(.A1(new_n761), .A2(new_n381), .B1(new_n763), .B2(new_n376), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G68), .B2(new_n795), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G97), .A2(new_n780), .B1(new_n777), .B2(G116), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1200), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n787), .A2(new_n1143), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n780), .A2(G132), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G128), .A2(new_n762), .B1(new_n764), .B2(G137), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n795), .A2(G150), .B1(G125), .B2(new_n777), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT114), .Z(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n266), .B(new_n245), .C1(new_n757), .C2(new_n771), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G124), .B2(new_n800), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT59), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1211), .B1(new_n1210), .B2(new_n1209), .C1(new_n1219), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n753), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n748), .B1(new_n202), .B2(new_n850), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1198), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1191), .B2(new_n745), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1197), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1128), .A2(new_n973), .A3(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n786), .A2(new_n296), .B1(new_n272), .B2(new_n770), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT121), .Z(new_n1234));
  OAI22_X1  g1034(.A1(new_n778), .A2(new_n520), .B1(new_n763), .B2(new_n381), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G116), .B2(new_n780), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT119), .Z(new_n1237));
  OAI21_X1  g1037(.A(new_n383), .B1(new_n757), .B2(new_n340), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1035), .B(new_n1239), .C1(G283), .C2(new_n762), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1234), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT122), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n787), .A2(G159), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n383), .B(new_n1202), .C1(G50), .C2(new_n795), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1143), .A2(new_n780), .B1(G132), .B2(new_n777), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n763), .A2(new_n838), .B1(new_n770), .B2(new_n1145), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G137), .B2(new_n762), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n753), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n749), .C1(G68), .C2(new_n1133), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n907), .B2(new_n804), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1125), .B2(new_n745), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1232), .A2(new_n1255), .ZN(G381));
  OR2_X1    g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1257), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1258), .ZN(G407));
  NAND2_X1  g1059(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT110), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1122), .A2(new_n1128), .A3(KEYINPUT110), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1260), .B1(new_n1265), .B2(new_n1121), .ZN(new_n1266));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G378), .B(new_n1229), .C1(new_n1193), .C2(new_n1196), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1228), .B1(new_n1194), .B2(new_n745), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1190), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1185), .A2(new_n1188), .A3(KEYINPUT118), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1192), .A3(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1276), .B2(new_n972), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1266), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1268), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT124), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G384), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n1106), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT123), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1231), .A2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1107), .A2(new_n712), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1284), .A2(new_n1285), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n828), .A2(KEYINPUT124), .A3(new_n852), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1290), .A2(new_n1255), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1281), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1289), .A2(new_n1291), .A3(new_n1281), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(G2897), .A3(new_n1268), .A4(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1289), .A2(new_n1291), .A3(new_n1281), .ZN(new_n1296));
  INV_X1    g1096(.A(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1268), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n1296), .A2(new_n1292), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1271), .B1(new_n1279), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT127), .B(new_n1271), .C1(new_n1279), .C2(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1279), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT62), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1279), .A2(new_n1308), .A3(new_n1305), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1303), .A2(new_n1304), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G390), .B(new_n1012), .C1(new_n1019), .C2(new_n971), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(G396), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(G390), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1014), .A2(new_n1020), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT126), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1014), .A2(new_n1020), .A3(new_n1317), .A4(new_n1314), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1313), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1314), .B1(new_n987), .B2(new_n1013), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1312), .B1(new_n1320), .B2(new_n1311), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1310), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1271), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1279), .A2(new_n1305), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(KEYINPUT63), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1306), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1279), .A2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1299), .B(new_n1295), .C1(new_n1279), .C2(new_n1329), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1326), .B(new_n1328), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(G405));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1266), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1305), .B1(new_n1334), .B2(new_n1272), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G378), .B1(new_n1197), .B2(new_n1229), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1272), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1296), .A2(new_n1292), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1335), .A2(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1322), .ZN(G402));
endmodule


