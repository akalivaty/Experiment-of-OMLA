//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n190), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n194), .A3(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT65), .B1(new_n191), .B2(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G143), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT82), .B1(new_n198), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n200), .B1(new_n203), .B2(G146), .ZN(new_n209));
  AND4_X1   g023(.A1(new_n204), .A2(new_n192), .A3(new_n194), .A4(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n192), .B2(new_n194), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(G128), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT82), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n202), .A4(new_n205), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n219), .A2(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .A4(new_n220), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n217), .A2(new_n218), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n196), .A2(G143), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n213), .B1(G143), .B2(new_n196), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n212), .A2(new_n233), .B1(new_n190), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n211), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT10), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT11), .A2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT11), .A4(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(G134), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT66), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT66), .B(new_n249), .C1(new_n246), .C2(G137), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n245), .B(new_n247), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT68), .A2(G131), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n249), .B1(new_n246), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n259), .A2(new_n251), .B1(new_n241), .B2(new_n244), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n247), .A3(new_n254), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n224), .A2(new_n227), .A3(new_n220), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT80), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n265), .A2(new_n269), .A3(new_n266), .A4(G101), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(G101), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n209), .B2(new_n210), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n212), .B2(new_n233), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n264), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n233), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n197), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n206), .A2(new_n274), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(new_n270), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT81), .A4(new_n273), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n239), .A2(new_n263), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G110), .B(G140), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT79), .ZN(new_n289));
  OR2_X1    g103(.A1(KEYINPUT71), .A2(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT71), .A2(G953), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G227), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n289), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n236), .A2(new_n231), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n217), .B2(new_n231), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n262), .A2(KEYINPUT83), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT12), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  INV_X1    g115(.A(new_n299), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n214), .A2(new_n202), .A3(new_n205), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n303), .A2(KEYINPUT82), .B1(new_n206), .B2(new_n208), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n230), .B1(new_n304), .B2(new_n216), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n301), .B(new_n302), .C1(new_n305), .C2(new_n297), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n239), .A2(new_n286), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT85), .B1(new_n309), .B2(new_n262), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n232), .A2(new_n238), .B1(new_n280), .B2(new_n285), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT85), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(new_n263), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n287), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n314), .B2(new_n294), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n315), .A2(G469), .A3(G902), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n312), .B1(new_n311), .B2(new_n263), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n309), .A2(KEYINPUT85), .A3(new_n262), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n296), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n239), .A2(new_n263), .A3(new_n286), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n307), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n287), .A2(KEYINPUT84), .A3(new_n300), .A4(new_n306), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n319), .B1(new_n324), .B2(new_n294), .ZN(new_n325));
  OAI21_X1  g139(.A(G469), .B1(new_n325), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n316), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT86), .B(G469), .C1(new_n325), .C2(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n189), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G137), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT77), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n292), .A2(G221), .A3(G234), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n334), .B(KEYINPUT78), .Z(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(G146), .B(new_n338), .C1(new_n342), .C2(new_n336), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  INV_X1    g158(.A(G119), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G110), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n190), .A2(G119), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT24), .B(G110), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT76), .B1(new_n351), .B2(new_n355), .ZN(new_n357));
  OAI221_X1 g171(.A(new_n343), .B1(G146), .B2(new_n342), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n338), .B1(new_n342), .B2(new_n336), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n196), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n343), .ZN(new_n361));
  OAI221_X1 g175(.A(new_n361), .B1(new_n350), .B2(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n335), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n334), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT25), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G217), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(G234), .B2(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(G902), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n364), .A2(new_n366), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT74), .ZN(new_n379));
  AOI21_X1  g193(.A(G131), .B1(new_n246), .B2(G137), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n245), .B(new_n380), .C1(new_n250), .C2(new_n252), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n247), .A2(KEYINPUT69), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n246), .A3(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n248), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT70), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(KEYINPUT70), .A3(new_n386), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n236), .ZN(new_n391));
  XOR2_X1   g205(.A(G116), .B(G119), .Z(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT2), .B(G113), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n262), .A2(new_n283), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n292), .A2(G210), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT27), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n292), .A2(new_n401), .A3(G210), .A4(new_n398), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G101), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n400), .B2(new_n402), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n236), .A2(new_n381), .A3(new_n386), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n387), .A2(new_n388), .B1(new_n211), .B2(new_n235), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n411), .A2(new_n390), .B1(new_n262), .B2(new_n283), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n412), .B2(new_n409), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n413), .B2(new_n394), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT31), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n395), .B1(new_n396), .B2(new_n408), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n397), .A2(KEYINPUT28), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n391), .A2(new_n396), .A3(new_n418), .A4(new_n395), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n414), .A2(new_n415), .B1(new_n420), .B2(new_n406), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n422));
  INV_X1    g236(.A(new_n410), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n409), .B1(new_n391), .B2(new_n396), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n394), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n407), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n422), .B1(new_n427), .B2(KEYINPUT31), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n415), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n421), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G472), .A2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT73), .Z(new_n432));
  OAI21_X1  g246(.A(new_n379), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n434));
  INV_X1    g248(.A(new_n432), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT72), .B1(new_n414), .B2(new_n415), .ZN(new_n436));
  AND4_X1   g250(.A1(KEYINPUT72), .A2(new_n425), .A3(new_n415), .A4(new_n426), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT74), .B(new_n435), .C1(new_n438), .C2(new_n421), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n429), .ZN(new_n441));
  INV_X1    g255(.A(new_n421), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n420), .A2(new_n406), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n445));
  INV_X1    g259(.A(new_n397), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n413), .B2(new_n394), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n444), .B(new_n445), .C1(new_n406), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n417), .A2(new_n419), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n395), .B2(new_n412), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n406), .A2(KEYINPUT29), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT75), .B(new_n367), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n395), .B1(new_n391), .B2(new_n396), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n454), .B(new_n451), .C1(new_n417), .C2(new_n419), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(G902), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n443), .A2(KEYINPUT32), .B1(new_n457), .B2(G472), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n378), .B1(new_n440), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT8), .Z(new_n462));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n392), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n345), .A3(G116), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G113), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n392), .A2(new_n393), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n462), .B1(new_n469), .B2(new_n230), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n464), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(KEYINPUT90), .A3(G113), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n470), .B1(new_n474), .B2(new_n230), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n283), .A2(G125), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n236), .A2(new_n340), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n478));
  INV_X1    g292(.A(G953), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G224), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n394), .A2(new_n273), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT88), .B1(new_n271), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n284), .A2(new_n490), .A3(new_n394), .A4(new_n273), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n469), .A2(new_n231), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(new_n461), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n461), .B(KEYINPUT89), .ZN(new_n496));
  AOI22_X1  g310(.A1(KEYINPUT6), .A2(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n485), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n460), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n499), .A3(new_n460), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G952), .ZN(new_n507));
  AOI211_X1 g321(.A(G953), .B(new_n507), .C1(G234), .C2(G237), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n367), .B(new_n292), .C1(G234), .C2(G237), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G116), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n226), .B1(new_n513), .B2(KEYINPUT14), .ZN(new_n514));
  XNOR2_X1  g328(.A(G116), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n192), .A2(new_n194), .A3(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n190), .A2(G143), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n246), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n246), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n515), .B(new_n226), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n517), .A2(new_n524), .A3(new_n518), .ZN(new_n525));
  OAI21_X1  g339(.A(G134), .B1(new_n517), .B2(new_n524), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n523), .B(new_n519), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n187), .A2(new_n373), .A3(G953), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n522), .A2(new_n527), .A3(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(KEYINPUT94), .A3(new_n530), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n367), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(G478), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(G478), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n367), .A3(new_n535), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n342), .B(G146), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n292), .A2(G143), .A3(G214), .A4(new_n398), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n290), .A2(G214), .A3(new_n398), .A4(new_n291), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n203), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n547));
  INV_X1    g361(.A(G131), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n542), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n547), .B(new_n548), .C1(new_n543), .C2(new_n545), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n342), .B(KEYINPUT19), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n548), .A3(new_n545), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n548), .B1(new_n543), .B2(new_n545), .ZN(new_n557));
  OAI221_X1 g371(.A(new_n343), .B1(G146), .B2(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G113), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n219), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n361), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n360), .A2(KEYINPUT91), .A3(new_n343), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OR3_X1    g382(.A1(new_n556), .A2(KEYINPUT17), .A3(new_n557), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n552), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n562), .B(new_n563), .C1(new_n570), .C2(new_n561), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT20), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n556), .A2(KEYINPUT17), .A3(new_n557), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n553), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n560), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n562), .A4(new_n563), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n560), .A2(KEYINPUT92), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n553), .B(new_n579), .C1(new_n573), .C2(new_n574), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n367), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n572), .A2(new_n578), .B1(new_n583), .B2(G475), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR4_X1   g399(.A1(new_n506), .A2(new_n511), .A3(new_n541), .A4(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n330), .A2(new_n459), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(new_n433), .A2(new_n439), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n441), .A2(new_n442), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n367), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n589), .A2(new_n378), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n330), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n504), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n501), .B2(new_n502), .ZN(new_n596));
  INV_X1    g410(.A(new_n511), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n528), .A2(KEYINPUT95), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n530), .A2(KEYINPUT96), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n533), .B2(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n599), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n534), .A2(new_n601), .A3(new_n535), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n367), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n536), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n584), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n596), .A2(new_n597), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n594), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND2_X1  g429(.A1(new_n503), .A2(new_n504), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n584), .A2(new_n541), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(new_n511), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT98), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  OR2_X1    g437(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n365), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n376), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n375), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n589), .A2(new_n628), .A3(new_n592), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n330), .A2(new_n586), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  AOI21_X1  g446(.A(new_n628), .B1(new_n440), .B2(new_n458), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n508), .B1(new_n509), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n616), .A2(new_n617), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n330), .A2(new_n633), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  XOR2_X1   g453(.A(new_n635), .B(KEYINPUT39), .Z(new_n640));
  NAND2_X1  g454(.A1(new_n330), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n503), .B(KEYINPUT38), .Z(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n443), .ZN(new_n646));
  INV_X1    g460(.A(new_n406), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n446), .B2(new_n454), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n427), .B2(new_n648), .ZN(new_n649));
  OAI221_X1 g463(.A(new_n440), .B1(new_n434), .B2(new_n646), .C1(new_n590), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n541), .A2(new_n504), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n584), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n628), .A2(new_n645), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n642), .A2(new_n643), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n195), .ZN(G45));
  NAND2_X1  g469(.A1(new_n611), .A2(new_n636), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT99), .B1(new_n616), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n610), .A2(new_n584), .A3(new_n635), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n596), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n330), .A2(new_n633), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  OAI21_X1  g476(.A(G469), .B1(new_n315), .B2(G902), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n321), .B1(new_n318), .B2(new_n317), .ZN(new_n664));
  OAI22_X1  g478(.A1(new_n664), .A2(new_n295), .B1(new_n307), .B2(new_n296), .ZN(new_n665));
  INV_X1    g479(.A(G469), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n367), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n663), .A2(new_n188), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n188), .A4(new_n667), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n459), .A2(new_n612), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  AND2_X1   g488(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(KEYINPUT101), .A3(new_n459), .A4(new_n618), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n459), .A2(new_n618), .A3(new_n670), .A4(new_n671), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  NAND2_X1  g495(.A1(new_n440), .A2(new_n458), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n585), .A2(new_n541), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n597), .A3(new_n683), .A4(new_n627), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n670), .A2(new_n596), .A3(new_n671), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n345), .ZN(G21));
  AOI22_X1  g501(.A1(new_n450), .A2(new_n647), .B1(new_n427), .B2(KEYINPUT31), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n432), .B1(new_n441), .B2(new_n688), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n592), .A2(new_n378), .A3(new_n511), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n502), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n652), .B1(new_n691), .B2(new_n500), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n503), .A2(KEYINPUT102), .A3(new_n652), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n696), .A3(new_n670), .A4(new_n671), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  INV_X1    g512(.A(new_n685), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n628), .A2(new_n592), .A3(new_n656), .A4(new_n689), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  NAND3_X1  g516(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n501), .A2(new_n705), .A3(new_n502), .A4(new_n504), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n189), .B1(new_n326), .B2(new_n667), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n659), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n434), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n443), .B2(KEYINPUT32), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n458), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n378), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT42), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n656), .A2(KEYINPUT42), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n459), .A2(new_n707), .A3(new_n708), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n548), .ZN(G33));
  NOR2_X1   g534(.A1(new_n617), .A2(new_n635), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n459), .A2(new_n707), .A3(new_n708), .A4(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n246), .ZN(G36));
  NAND2_X1  g539(.A1(G469), .A2(G902), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n325), .A2(KEYINPUT45), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n666), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n325), .A2(KEYINPUT45), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n727), .B(new_n729), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n730), .B(KEYINPUT106), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n727), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n726), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n316), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n729), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n733), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT108), .A3(KEYINPUT46), .A4(new_n726), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT46), .B(new_n726), .C1(new_n734), .C2(new_n736), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n188), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n627), .B1(new_n589), .B2(new_n592), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(KEYINPUT109), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(KEYINPUT109), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n585), .A2(new_n610), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT43), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n707), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT44), .B1(new_n753), .B2(new_n755), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n749), .A2(new_n760), .A3(new_n640), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n748), .B(new_n763), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n758), .A2(new_n682), .A3(new_n714), .A4(new_n656), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  NAND3_X1  g581(.A1(new_n714), .A2(new_n188), .A3(new_n505), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT110), .Z(new_n769));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n663), .A2(new_n667), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n769), .B(new_n754), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT111), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n650), .B(new_n645), .C1(new_n770), .C2(new_n772), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n330), .B(new_n586), .C1(new_n459), .C2(new_n629), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n704), .A2(new_n683), .A3(new_n706), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n330), .A2(new_n633), .A3(new_n636), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n611), .B1(new_n541), .B2(new_n584), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n506), .A3(new_n511), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n330), .A2(new_n593), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n700), .A2(new_n707), .A3(new_n708), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n778), .A2(new_n780), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n724), .A2(new_n785), .A3(new_n719), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n672), .A2(new_n697), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n686), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n680), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n680), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n790), .A3(KEYINPUT113), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n635), .B1(new_n694), .B2(new_n695), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n650), .A2(new_n794), .A3(new_n628), .A4(new_n708), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n701), .A2(new_n638), .A3(new_n661), .A4(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT52), .Z(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n788), .A2(new_n680), .A3(new_n791), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n791), .B1(new_n788), .B2(new_n680), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n801), .B2(new_n786), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n777), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n786), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n796), .B(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n788), .A2(new_n680), .A3(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n803), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n777), .C1(new_n798), .C2(new_n802), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n798), .A2(new_n802), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n810), .B1(new_n816), .B2(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n592), .A2(new_n689), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n714), .A2(new_n755), .A3(new_n508), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n707), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n748), .B(KEYINPUT47), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n771), .B(KEYINPUT116), .Z(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n188), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT117), .Z(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n675), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n758), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n508), .A3(new_n755), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n819), .A2(new_n627), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n714), .A2(new_n508), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n827), .A2(new_n650), .A3(new_n758), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n585), .A2(new_n609), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n675), .A3(new_n595), .A4(new_n644), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n818), .B1(new_n826), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n829), .A2(new_n715), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT48), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n845), .A2(KEYINPUT120), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n833), .A2(new_n611), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n507), .B(G953), .C1(new_n820), .C2(new_n699), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n850));
  OAI211_X1 g664(.A(new_n848), .B(new_n849), .C1(new_n845), .C2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n707), .B(new_n820), .C1(new_n764), .C2(new_n824), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n835), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n847), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n817), .A2(new_n842), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(G952), .A2(G953), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n776), .B1(new_n855), .B2(new_n856), .ZN(G75));
  AOI21_X1  g671(.A(new_n367), .B1(new_n803), .B2(new_n808), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT56), .B1(new_n858), .B2(G210), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n497), .A2(new_n498), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n485), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n292), .A2(G952), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n859), .A2(KEYINPUT121), .A3(new_n862), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n859), .B2(new_n862), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(G51));
  XOR2_X1   g683(.A(new_n726), .B(KEYINPUT57), .Z(new_n870));
  AOI21_X1  g684(.A(new_n809), .B1(new_n803), .B2(new_n808), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n810), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n665), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n858), .A2(new_n733), .A3(new_n741), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n864), .B1(new_n873), .B2(new_n874), .ZN(G54));
  NAND2_X1  g689(.A1(new_n576), .A2(new_n562), .ZN(new_n876));
  INV_X1    g690(.A(new_n858), .ZN(new_n877));
  NAND2_X1  g691(.A1(KEYINPUT58), .A2(G475), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n865), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n877), .A2(new_n876), .A3(new_n878), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(G60));
  NAND2_X1  g696(.A1(new_n604), .A2(new_n605), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n884));
  NAND2_X1  g698(.A1(G478), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n817), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n883), .A2(new_n886), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n803), .A2(new_n808), .ZN(new_n891));
  INV_X1    g705(.A(new_n809), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n803), .A2(new_n808), .A3(new_n809), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n888), .B1(new_n895), .B2(new_n864), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n889), .B1(new_n810), .B2(new_n871), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT123), .A3(new_n865), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n887), .A2(new_n896), .A3(new_n898), .ZN(G63));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n364), .A2(new_n366), .ZN(new_n901));
  INV_X1    g715(.A(new_n891), .ZN(new_n902));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n865), .ZN(new_n906));
  INV_X1    g720(.A(new_n625), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n902), .A2(new_n907), .A3(new_n904), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n900), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n908), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n865), .A4(new_n905), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(G66));
  INV_X1    g726(.A(new_n510), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n479), .B1(new_n913), .B2(G224), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n801), .A2(new_n783), .A3(new_n778), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n292), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n860), .B1(G898), .B2(new_n292), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT124), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(G69));
  INV_X1    g733(.A(new_n292), .ZN(new_n920));
  INV_X1    g734(.A(G227), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n634), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n413), .B(new_n554), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n634), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n715), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n749), .A2(new_n640), .A3(new_n696), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n701), .A2(new_n638), .A3(new_n661), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n724), .A2(new_n932), .A3(new_n719), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n766), .A2(new_n761), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n934), .B2(new_n292), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n926), .A2(new_n920), .ZN(new_n936));
  INV_X1    g750(.A(new_n765), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n822), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n654), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT62), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n758), .A2(new_n781), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n459), .A3(new_n330), .A4(new_n640), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n761), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n924), .B(new_n925), .C1(new_n935), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n931), .A2(new_n761), .A3(new_n933), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n926), .B(new_n928), .C1(new_n949), .C2(new_n920), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(new_n945), .A3(new_n923), .A4(new_n922), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n947), .A2(new_n951), .ZN(G72));
  XOR2_X1   g766(.A(new_n447), .B(KEYINPUT127), .Z(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n647), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n938), .A2(new_n948), .A3(new_n915), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT63), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n953), .A2(new_n647), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n938), .A2(new_n944), .A3(new_n915), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n957), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n961), .A3(new_n865), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n447), .A2(new_n406), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n957), .B1(new_n963), .B2(new_n427), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n816), .B2(new_n964), .ZN(G57));
endmodule


