//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G68), .A2(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n208), .B1(new_n202), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g0010(.A1(G77), .A2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n210), .B(new_n211), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n218), .B1(new_n217), .B2(new_n216), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n224), .B(new_n227), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n220), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n209), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n219), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT8), .A2(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT68), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n229), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n203), .A2(KEYINPUT70), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT69), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n268), .B1(new_n262), .B2(new_n264), .C1(new_n260), .C2(new_n261), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n229), .B1(new_n201), .B2(new_n202), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n266), .A2(new_n267), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n228), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n255), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n253), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n202), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT9), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n228), .ZN(new_n286));
  AND2_X1   g0086(.A1(G1), .A2(G13), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n283), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G226), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n286), .B2(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1698), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(G222), .B1(new_n300), .B2(G77), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT3), .B(G33), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G223), .A3(G1698), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n285), .A2(new_n228), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n291), .B(new_n294), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT67), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n308), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G190), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n307), .B(KEYINPUT67), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n277), .A2(new_n202), .ZN(new_n315));
  AOI211_X1 g0115(.A(new_n255), .B(new_n315), .C1(new_n272), .C2(new_n274), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT9), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n280), .A2(new_n312), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n319));
  AOI22_X1  g0119(.A1(G200), .A2(new_n313), .B1(new_n316), .B2(KEYINPUT9), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n312), .A4(new_n280), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n311), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n302), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n302), .A2(G232), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n330), .B1(new_n332), .B2(new_n209), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n305), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n290), .A2(G238), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n294), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n337), .B(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT14), .B1(new_n339), .B2(new_n326), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(G179), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n337), .B(KEYINPUT13), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(G169), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n347), .B1(new_n261), .B2(new_n348), .C1(new_n264), .C2(new_n202), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(new_n274), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(KEYINPUT11), .B1(G68), .B2(new_n276), .ZN(new_n351));
  INV_X1    g0151(.A(new_n254), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n346), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n354), .C1(KEYINPUT11), .C2(new_n350), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT73), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n274), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n232), .B1(new_n258), .B2(new_n346), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n300), .B2(new_n229), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n298), .A2(new_n299), .A3(new_n362), .A4(G20), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n358), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n298), .A2(new_n299), .A3(G20), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT74), .B1(new_n368), .B2(KEYINPUT7), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n295), .A2(new_n229), .A3(new_n296), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n362), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n363), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT16), .B(new_n360), .C1(new_n373), .C2(new_n346), .ZN(new_n374));
  INV_X1    g0174(.A(new_n260), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n277), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n260), .A2(new_n254), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n367), .A2(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(G226), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n379));
  OAI211_X1 g0179(.A(G223), .B(new_n331), .C1(new_n298), .C2(new_n299), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n305), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n290), .A2(G232), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n294), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT75), .B1(new_n385), .B2(G190), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n382), .A2(new_n305), .B1(new_n293), .B2(new_n283), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT75), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .A4(new_n384), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n378), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n378), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n367), .A2(new_n374), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n376), .A2(new_n377), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n385), .A2(new_n324), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n326), .B1(new_n389), .B2(new_n384), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT18), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n356), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n339), .A2(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n342), .A2(G200), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G20), .A2(G77), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n263), .B(KEYINPUT71), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT8), .B(G58), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT15), .B(G87), .Z(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n416), .B1(new_n417), .B2(new_n418), .C1(new_n261), .C2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n274), .B1(new_n348), .B2(new_n352), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n276), .A2(G77), .ZN(new_n423));
  XOR2_X1   g0223(.A(new_n423), .B(KEYINPUT72), .Z(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n302), .A2(G238), .A3(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G107), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n426), .B1(new_n427), .B2(new_n302), .C1(new_n333), .C2(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n305), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n290), .A2(G244), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n294), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n425), .B1(G179), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n431), .A2(new_n326), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n357), .A2(new_n411), .A3(new_n415), .A4(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n425), .B1(G200), .B2(new_n431), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n431), .A2(new_n391), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n329), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT21), .ZN(new_n442));
  OAI211_X1 g0242(.A(G264), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n302), .A2(KEYINPUT78), .A3(G264), .A4(G1698), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G303), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n332), .A2(new_n215), .B1(new_n448), .B2(new_n302), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n305), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n253), .A2(G45), .ZN(new_n452));
  OR2_X1    g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n286), .B2(new_n289), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G270), .B1(new_n293), .B2(new_n455), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n450), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT81), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n254), .B2(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n253), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n254), .A2(new_n464), .A3(new_n228), .A4(new_n273), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(new_n219), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n273), .A2(new_n228), .B1(G20), .B2(new_n219), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n229), .C1(G33), .C2(new_n214), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n465), .A2(KEYINPUT80), .A3(new_n219), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n473), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(KEYINPUT81), .A3(new_n466), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G169), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n442), .B1(new_n460), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n450), .A2(new_n457), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT79), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(KEYINPUT21), .A3(G169), .A4(new_n480), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n483), .A2(new_n324), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n480), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n482), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n387), .B1(new_n484), .B2(new_n485), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT82), .B1(new_n491), .B2(new_n480), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(new_n480), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n460), .C2(new_n387), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n460), .A2(G190), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT83), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n490), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n254), .A2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n465), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G97), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n361), .B2(new_n363), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n214), .A2(new_n427), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n205), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n427), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G20), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n264), .A2(new_n348), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT76), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n516), .A3(new_n274), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n515), .B2(new_n274), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n503), .B(new_n505), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(new_n331), .C1(new_n298), .C2(new_n299), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n302), .A2(KEYINPUT4), .A3(G244), .A4(new_n331), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n302), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n468), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n305), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n293), .A2(new_n455), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n456), .A2(G257), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n324), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n525), .A2(new_n305), .B1(new_n293), .B2(new_n455), .ZN(new_n530));
  AOI21_X1  g0330(.A(G169), .B1(new_n530), .B2(new_n528), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n370), .A2(new_n362), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n300), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n427), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n229), .B1(new_n509), .B2(new_n510), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n536), .A2(new_n537), .A3(new_n513), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT76), .B1(new_n538), .B2(new_n358), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n515), .A2(new_n516), .A3(new_n274), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n502), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n530), .A2(new_n391), .A3(new_n528), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(G200), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n544), .A3(new_n505), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n465), .A2(new_n427), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT22), .B(G87), .C1(new_n298), .C2(new_n299), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n229), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n302), .A2(new_n229), .A3(G87), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI211_X1 g0354(.A(G20), .B(new_n427), .C1(new_n554), .C2(KEYINPUT84), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(KEYINPUT84), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT24), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n549), .A2(new_n229), .B1(new_n551), .B2(new_n552), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n557), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n546), .B1(new_n563), .B2(new_n274), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n302), .A2(G257), .A3(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n302), .A2(KEYINPUT85), .A3(G257), .A4(G1698), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n297), .A2(G250), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n305), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n456), .A2(G264), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(G190), .A3(new_n527), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n527), .A3(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n254), .A2(G107), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT25), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n564), .A2(new_n574), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n533), .A2(new_n545), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n297), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n302), .A2(G244), .A3(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n305), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n285), .A2(new_n284), .A3(new_n228), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT66), .B1(new_n287), .B2(new_n288), .ZN(new_n586));
  OAI211_X1 g0386(.A(G250), .B(new_n452), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n284), .A2(new_n253), .A3(G45), .A4(G274), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n587), .A2(KEYINPUT77), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT77), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n584), .B(G190), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n419), .A2(new_n254), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n229), .B1(new_n330), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n205), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n594), .A2(new_n596), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n302), .A2(new_n229), .A3(G68), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n358), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n592), .B(new_n600), .C1(G87), .C2(new_n504), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n306), .B1(new_n581), .B2(new_n582), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n587), .A2(new_n588), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT77), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n587), .A2(KEYINPUT77), .A3(new_n588), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n591), .B(new_n601), .C1(new_n607), .C2(new_n387), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n584), .B(new_n324), .C1(new_n589), .C2(new_n590), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n600), .A2(new_n592), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n420), .B2(new_n465), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n611), .C1(new_n607), .C2(G169), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n558), .A2(KEYINPUT24), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n561), .B1(new_n560), .B2(new_n557), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n274), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n546), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n578), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n575), .A2(G179), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n575), .A2(new_n326), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n580), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n441), .A2(new_n501), .A3(new_n622), .ZN(G372));
  NAND3_X1  g0423(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n326), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n530), .A2(new_n324), .A3(new_n528), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n541), .B2(new_n505), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n607), .B2(new_n387), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n610), .B1(new_n595), .B2(new_n465), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n607), .B2(G190), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT86), .A3(G200), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n628), .A2(new_n629), .A3(new_n612), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n519), .A2(new_n532), .A3(new_n608), .A4(new_n612), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n637), .A2(new_n612), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n533), .A2(new_n545), .A3(new_n579), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n482), .A3(new_n487), .A4(new_n489), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n612), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n441), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n328), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n401), .B2(new_n405), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n378), .A2(new_n404), .A3(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n408), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n401), .A2(new_n405), .A3(new_n650), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT87), .B1(new_n378), .B2(new_n404), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n356), .A2(new_n345), .B1(new_n415), .B2(new_n434), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n398), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n649), .B1(new_n659), .B2(new_n323), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n648), .A2(new_n660), .ZN(G369));
  INV_X1    g0461(.A(G13), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G20), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n253), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n253), .A2(new_n229), .A3(G13), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n667), .A3(G213), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n494), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n501), .B(new_n490), .S(new_n674), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n618), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n621), .B1(new_n579), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n642), .A2(new_n672), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(G330), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n490), .A2(new_n673), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(new_n681), .A3(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n225), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n596), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n233), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n482), .A2(new_n487), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n489), .A4(new_n642), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n580), .A2(new_n644), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n643), .A2(KEYINPUT90), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n699));
  INV_X1    g0499(.A(new_n612), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n645), .A2(new_n628), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(KEYINPUT26), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT91), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n672), .B1(new_n640), .B2(new_n646), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n703), .A2(new_n708), .A3(KEYINPUT29), .A4(new_n673), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n498), .A2(new_n500), .ZN(new_n711));
  INV_X1    g0511(.A(new_n490), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n622), .A4(new_n673), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n572), .A2(new_n573), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n634), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n488), .A3(new_n543), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n488), .A4(new_n543), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n543), .A2(new_n607), .A3(G179), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n721), .A2(new_n486), .A3(new_n575), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n672), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n725), .B(new_n672), .C1(new_n720), .C2(new_n722), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n713), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n710), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n692), .B1(new_n731), .B2(G1), .ZN(G364));
  AOI21_X1  g0532(.A(new_n253), .B1(new_n663), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n687), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n248), .A2(G45), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n686), .A2(new_n302), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(G45), .C2(new_n233), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n302), .A2(new_n225), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n738), .B1(G116), .B2(new_n225), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT92), .B1(G13), .B2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(KEYINPUT92), .A2(G13), .A3(G33), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n228), .B1(G20), .B2(new_n326), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n229), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G159), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT32), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n229), .B1(new_n751), .B2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n755), .B1(G97), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n302), .B1(new_n761), .B2(new_n346), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n324), .A2(G200), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(new_n750), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n387), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n348), .B1(new_n427), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n229), .A2(new_n391), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n766), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n762), .B(new_n768), .C1(G87), .C2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n759), .A2(new_n391), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT93), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n769), .A2(new_n763), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n773), .B1(new_n202), .B2(new_n778), .C1(new_n258), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n761), .B1(KEYINPUT33), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(KEYINPUT33), .B2(new_n781), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n300), .C1(new_n784), .C2(new_n756), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G311), .B2(new_n764), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(G303), .ZN(new_n787));
  INV_X1    g0587(.A(new_n778), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G326), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n779), .A2(new_n790), .B1(new_n767), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n752), .B(KEYINPUT94), .Z(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(G329), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n786), .A2(new_n787), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n780), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n747), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n735), .B(new_n749), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  INV_X1    g0602(.A(new_n746), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n802), .C1(new_n675), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n675), .A2(G330), .ZN(new_n805));
  INV_X1    g0605(.A(new_n735), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n675), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(G396));
  INV_X1    g0609(.A(KEYINPUT98), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n435), .A2(new_n672), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n672), .A2(new_n425), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n439), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n435), .B2(new_n813), .ZN(new_n814));
  AND4_X1   g0614(.A1(new_n810), .A2(new_n647), .A3(new_n673), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n810), .B1(new_n706), .B2(new_n814), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n816), .B1(new_n706), .B2(new_n814), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n729), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n735), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n300), .B1(new_n770), .B2(new_n427), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n767), .A2(new_n595), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n794), .C2(G311), .ZN(new_n822));
  INV_X1    g0622(.A(new_n779), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(G294), .B1(new_n757), .B2(G97), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n448), .C2(new_n778), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n764), .A2(G116), .B1(new_n760), .B2(G283), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT97), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n770), .A2(new_n202), .B1(new_n756), .B2(new_n258), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n764), .A2(G159), .B1(new_n760), .B2(G150), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n779), .C1(new_n778), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT34), .Z(new_n834));
  INV_X1    g0634(.A(new_n767), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n829), .B(new_n834), .C1(G68), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n300), .B1(new_n794), .B2(G132), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n745), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n747), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT96), .Z(new_n841));
  OAI22_X1  g0641(.A1(new_n838), .A2(new_n798), .B1(G77), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n814), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n806), .B(new_n842), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n819), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  OAI211_X1 g0646(.A(G116), .B(new_n230), .C1(new_n511), .C2(KEYINPUT35), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT36), .ZN(new_n851));
  INV_X1    g0651(.A(new_n258), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n348), .B(new_n233), .C1(G68), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n346), .A2(G50), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n662), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n851), .B1(new_n253), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  INV_X1    g0658(.A(KEYINPUT39), .ZN(new_n859));
  INV_X1    g0659(.A(new_n669), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n360), .B1(new_n373), .B2(new_n346), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n366), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n360), .B1(KEYINPUT102), .B2(KEYINPUT16), .C1(new_n373), .C2(new_n346), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n274), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n860), .B1(new_n865), .B2(new_n400), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n398), .B2(new_n410), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n865), .A2(new_n400), .B1(new_n404), .B2(new_n860), .ZN(new_n868));
  INV_X1    g0668(.A(new_n394), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n401), .A2(new_n669), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(new_n406), .A3(new_n872), .A4(new_n394), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n395), .A2(new_n397), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT18), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT18), .B1(new_n654), .B2(new_n655), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n871), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n651), .A2(new_n652), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n871), .A2(new_n394), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n879), .A2(new_n880), .B1(new_n883), .B2(new_n873), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n859), .B(new_n875), .C1(new_n884), .C2(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n883), .A2(new_n873), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n871), .B1(new_n657), .B2(new_n876), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n859), .A4(new_n875), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT103), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n870), .A2(new_n873), .ZN(new_n894));
  INV_X1    g0694(.A(new_n866), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n408), .B1(new_n401), .B2(new_n405), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n378), .A2(new_n404), .A3(KEYINPUT18), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n898), .B2(new_n876), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n888), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n875), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n893), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n902));
  AOI211_X1 g0702(.A(KEYINPUT103), .B(new_n859), .C1(new_n900), .C2(new_n875), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n887), .B(new_n892), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n357), .A2(new_n672), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n653), .A2(new_n656), .A3(new_n860), .ZN(new_n907));
  INV_X1    g0707(.A(new_n811), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n815), .B2(new_n816), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n357), .B(new_n415), .C1(new_n412), .C2(new_n673), .ZN(new_n910));
  INV_X1    g0710(.A(new_n415), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n356), .B(new_n672), .C1(new_n911), .C2(new_n345), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n901), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n906), .A2(new_n907), .A3(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n705), .A2(new_n441), .A3(new_n707), .A4(new_n709), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n660), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n843), .B1(new_n713), .B2(new_n727), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n901), .A3(new_n913), .ZN(new_n920));
  OR2_X1    g0720(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n921));
  NAND2_X1  g0721(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n891), .A2(new_n875), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(KEYINPUT40), .A3(new_n913), .A4(new_n919), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n441), .A2(new_n728), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G330), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n918), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n663), .A2(new_n253), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n858), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT106), .Z(G367));
  AOI22_X1  g0734(.A1(new_n764), .A2(G50), .B1(new_n760), .B2(G159), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT112), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n302), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n835), .A2(G77), .B1(new_n753), .B2(G137), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n262), .B2(new_n779), .C1(new_n258), .C2(new_n770), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n937), .B(new_n939), .C1(G68), .C2(new_n757), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(KEYINPUT112), .B2(new_n935), .C1(new_n831), .C2(new_n778), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n835), .A2(G97), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n942), .B1(new_n448), .B2(new_n779), .C1(new_n781), .C2(new_n752), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n770), .A2(new_n219), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT46), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n761), .A2(new_n784), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n300), .B1(new_n756), .B2(new_n427), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n943), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(G311), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n948), .B1(new_n791), .B2(new_n765), .C1(new_n949), .C2(new_n778), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n806), .B1(new_n952), .B2(new_n747), .ZN(new_n953));
  INV_X1    g0753(.A(new_n737), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n748), .B1(new_n225), .B2(new_n420), .C1(new_n240), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n672), .A2(new_n632), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n700), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n644), .B2(new_n956), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n953), .B(new_n955), .C1(new_n803), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n672), .A2(new_n519), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n545), .A3(new_n533), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n628), .A2(new_n672), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n533), .B1(new_n961), .B2(new_n642), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n673), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT42), .B1(new_n684), .B2(new_n964), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n958), .B(KEYINPUT107), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n965), .A2(new_n972), .A3(new_n967), .A4(new_n968), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT108), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n979), .A3(new_n975), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n680), .A2(new_n964), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n982), .A3(new_n980), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n963), .B(new_n681), .C1(new_n677), .C2(new_n682), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT110), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT110), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n681), .B1(new_n677), .B2(new_n682), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n964), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n993), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n680), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n992), .A2(new_n680), .A3(new_n993), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n679), .B(new_n682), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1004), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n805), .A2(KEYINPUT111), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n731), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n687), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n734), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n959), .B1(new_n986), .B2(new_n1013), .ZN(G387));
  NAND3_X1  g0814(.A1(new_n731), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n688), .B1(new_n1008), .B2(new_n730), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n679), .A2(new_n803), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n737), .B1(new_n244), .B2(new_n282), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n689), .B2(new_n740), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G116), .B(new_n596), .C1(G68), .C2(G77), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT50), .B1(new_n418), .B2(G50), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n418), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n282), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1020), .A2(new_n1024), .B1(new_n427), .B2(new_n686), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n748), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n735), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT113), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n764), .A2(G303), .B1(new_n760), .B2(G311), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n781), .B2(new_n779), .C1(new_n778), .C2(new_n790), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n791), .B2(new_n756), .C1(new_n784), .C2(new_n770), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n753), .A2(G326), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n302), .B1(new_n835), .B2(G116), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n420), .A2(new_n756), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n770), .A2(new_n348), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G150), .B2(new_n753), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n202), .B2(new_n779), .C1(new_n346), .C2(new_n765), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n375), .C2(new_n760), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n788), .A2(G159), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1043), .A2(new_n302), .A3(new_n942), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1028), .B1(new_n798), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1017), .B1(new_n733), .B2(new_n1008), .C1(new_n1018), .C2(new_n1048), .ZN(G393));
  NAND3_X1  g0849(.A1(new_n1000), .A2(new_n734), .A3(new_n1001), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n778), .A2(new_n781), .B1(new_n949), .B2(new_n779), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n770), .A2(new_n791), .B1(new_n752), .B2(new_n790), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n300), .B1(new_n761), .B2(new_n448), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n767), .A2(new_n427), .B1(new_n756), .B2(new_n219), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1052), .B(new_n1056), .C1(new_n784), .C2(new_n765), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n788), .A2(G150), .B1(G159), .B2(new_n823), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n756), .A2(new_n348), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n765), .A2(new_n418), .B1(new_n752), .B2(new_n831), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G68), .C2(new_n771), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n300), .B(new_n821), .C1(G50), .C2(new_n760), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n806), .B1(new_n1066), .B2(new_n747), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n748), .B1(new_n214), .B2(new_n225), .C1(new_n251), .C2(new_n954), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n963), .C2(new_n803), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1050), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1015), .A2(new_n1002), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n687), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1015), .A2(new_n1002), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(G390));
  AOI21_X1  g0875(.A(new_n905), .B1(new_n891), .B2(new_n875), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n813), .A2(new_n435), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n703), .A2(new_n673), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n908), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n913), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n905), .B1(new_n909), .B2(new_n913), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(new_n904), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n919), .A2(G330), .A3(new_n913), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1081), .B(KEYINPUT115), .C1(new_n1082), .C2(new_n904), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1086), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1083), .A2(new_n1084), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n913), .B1(new_n919), .B2(G330), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n909), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT116), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1079), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT116), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n909), .C1(new_n1086), .C2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G330), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n916), .B(new_n660), .C1(new_n1100), .C2(new_n927), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1091), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1088), .A2(new_n1090), .A3(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n687), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n904), .A2(new_n745), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n302), .B1(new_n765), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n770), .A2(new_n262), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n757), .A2(G159), .B1(new_n760), .B2(G137), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1111), .B(new_n1115), .C1(G125), .C2(new_n794), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  INV_X1    g0917(.A(G132), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n778), .A2(new_n1117), .B1(new_n1118), .B2(new_n779), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT117), .Z(new_n1120));
  OAI211_X1 g0920(.A(new_n1116), .B(new_n1120), .C1(new_n202), .C2(new_n767), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n765), .A2(new_n214), .B1(new_n346), .B2(new_n767), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n794), .B2(G294), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n300), .B1(new_n761), .B2(new_n427), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1060), .B(new_n1124), .C1(G87), .C2(new_n771), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n219), .B2(new_n779), .C1(new_n791), .C2(new_n778), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n798), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n841), .A2(new_n375), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1108), .A2(new_n806), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1091), .B2(new_n734), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1107), .A2(new_n1131), .ZN(G378));
  NOR2_X1   g0932(.A1(new_n316), .A2(new_n860), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n329), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT55), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1133), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n323), .A2(new_n328), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n323), .B2(new_n328), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1133), .B(new_n649), .C1(new_n319), .C2(new_n322), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT55), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT56), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT56), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n926), .B2(new_n1100), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT56), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n1142), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1148), .A2(G330), .A3(new_n923), .A4(new_n925), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n915), .A2(KEYINPUT119), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1146), .A2(new_n1149), .A3(new_n915), .A4(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1103), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n1101), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n915), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1150), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1146), .A2(new_n1149), .A3(new_n915), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1155), .B2(new_n1101), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n687), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1154), .A2(new_n734), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n761), .A2(new_n1118), .B1(new_n262), .B2(new_n756), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n765), .A2(new_n832), .B1(new_n1117), .B2(new_n779), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n788), .C2(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n770), .B2(new_n1110), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT59), .Z(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n753), .B2(G124), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G33), .B1(new_n835), .B2(G159), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G50), .B1(new_n296), .B2(new_n281), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n778), .A2(new_n219), .B1(new_n346), .B2(new_n756), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT118), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n852), .A2(new_n835), .B1(new_n764), .B2(new_n419), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n427), .B2(new_n779), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1040), .B(new_n1178), .C1(G283), .C2(new_n794), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G41), .B(new_n302), .C1(G97), .C2(new_n760), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1176), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT58), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1174), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1173), .B(new_n1183), .C1(new_n1182), .C2(new_n1181), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n841), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1184), .A2(new_n747), .B1(new_n202), .B2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n735), .B(new_n1186), .C1(new_n1145), .C2(new_n745), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1165), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n1189), .ZN(G375));
  NAND4_X1  g0990(.A1(new_n1101), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1103), .A2(new_n1012), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n793), .A2(new_n448), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n300), .B1(new_n761), .B2(new_n219), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n420), .A2(new_n756), .B1(new_n348), .B2(new_n767), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n214), .A2(new_n770), .B1(new_n779), .B2(new_n791), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n427), .B2(new_n765), .C1(new_n784), .C2(new_n778), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT120), .Z(new_n1199));
  NOR2_X1   g0999(.A1(new_n779), .A2(new_n832), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n756), .A2(new_n202), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n302), .B1(new_n767), .B2(new_n258), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G159), .C2(new_n771), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n1117), .B2(new_n793), .C1(new_n262), .C2(new_n765), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT121), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n788), .A2(G132), .B1(new_n760), .B2(new_n1109), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1199), .B1(new_n1200), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n735), .B1(new_n745), .B2(new_n913), .C1(new_n1211), .C2(new_n798), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n346), .B2(new_n1185), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1099), .B2(new_n734), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1192), .A2(new_n1214), .ZN(G381));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G387), .A2(G390), .A3(G384), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1164), .A2(new_n1217), .A3(new_n1189), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1214), .A3(new_n1192), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1219), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(new_n1225), .ZN(G407));
  INV_X1    g1026(.A(G213), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1105), .A2(new_n1102), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n688), .B1(new_n1228), .B2(new_n1162), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1188), .B1(new_n1229), .B2(new_n1158), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1217), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G343), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1227), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(G409));
  XOR2_X1   g1039(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1240));
  AND3_X1   g1040(.A1(new_n1107), .A2(new_n1131), .A3(new_n1187), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1012), .B(new_n1154), .C1(new_n1155), .C2(new_n1101), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n734), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1227), .A2(G343), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n1230), .C2(new_n1217), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1099), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(KEYINPUT60), .A4(new_n1101), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT125), .B1(new_n1191), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1191), .A2(new_n1253), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n688), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1257), .A2(G384), .A3(new_n1214), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1257), .B2(new_n1214), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G2897), .B(new_n1247), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1214), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n845), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(G384), .A3(new_n1214), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(G2897), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1240), .B1(new_n1249), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1247), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n1217), .C2(new_n1230), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT62), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1267), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1221), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1074), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n688), .B1(new_n1015), .B2(new_n1002), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1070), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G387), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1276), .B(new_n1277), .C1(new_n1281), .C2(KEYINPUT126), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G390), .B(new_n959), .C1(new_n1013), .C2(new_n986), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1280), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1282), .B(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1275), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1272), .B2(new_n1268), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1270), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1217), .B1(new_n1164), .B2(new_n1189), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1107), .A2(new_n1131), .A3(new_n1187), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1248), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1269), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1292), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1286), .B1(new_n1297), .B2(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1291), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(new_n1300), .ZN(G405));
  OR2_X1    g1101(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1302), .B(new_n1303), .C1(new_n1232), .C2(new_n1292), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1286), .A2(new_n1231), .A3(new_n1272), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1269), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1269), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(G402));
endmodule


