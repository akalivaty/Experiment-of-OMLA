//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(G197gat), .ZN(new_n205));
  INV_X1    g004(.A(G204gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  AND2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n207), .A2(new_n208), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n213));
  INV_X1    g012(.A(new_n211), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n210), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G226gat), .A2(G233gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT26), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(KEYINPUT27), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT28), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n229), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n233), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n247), .B1(KEYINPUT65), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n249), .A2(new_n251), .A3(new_n254), .A4(new_n250), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT25), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT25), .A4(new_n246), .ZN(new_n257));
  INV_X1    g056(.A(new_n250), .ZN(new_n258));
  AND2_X1   g057(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n233), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT24), .B1(new_n227), .B2(KEYINPUT66), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(KEYINPUT66), .B2(new_n227), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n257), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n242), .B1(new_n256), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n220), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n270));
  INV_X1    g069(.A(new_n247), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n255), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n265), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n242), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(KEYINPUT68), .B(new_n229), .C1(new_n237), .C2(new_n241), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n268), .A2(new_n269), .B1(new_n280), .B2(new_n220), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT29), .B1(new_n276), .B2(new_n242), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT78), .B1(new_n282), .B2(new_n220), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n218), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(new_n220), .ZN(new_n287));
  INV_X1    g086(.A(new_n239), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n235), .B1(new_n261), .B2(KEYINPUT27), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(KEYINPUT28), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n274), .A2(new_n275), .B1(new_n291), .B2(new_n229), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n280), .A2(new_n287), .B1(new_n292), .B2(new_n220), .ZN(new_n293));
  INV_X1    g092(.A(new_n218), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT30), .B(new_n204), .C1(new_n284), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT79), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n269), .B(new_n219), .C1(new_n292), .C2(KEYINPUT29), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n220), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n294), .ZN(new_n301));
  INV_X1    g100(.A(new_n295), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT30), .A4(new_n204), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n284), .A2(new_n295), .A3(new_n204), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n204), .B1(new_n284), .B2(new_n295), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G113gat), .A2(G120gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g112(.A1(G113gat), .A2(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  INV_X1    g120(.A(G127gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(G134gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n328));
  OAI21_X1  g127(.A(G120gat), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n313), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G155gat), .B(G162gat), .Z(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT80), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n332), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G148gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT81), .B1(new_n340), .B2(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(G141gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  OR2_X1    g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n326), .A2(new_n331), .A3(new_n339), .A4(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(G134gat), .A3(new_n316), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n323), .A3(new_n324), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n319), .A2(G127gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n322), .A2(G134gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G113gat), .B2(G120gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n356), .A2(new_n315), .B1(new_n362), .B2(new_n329), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n343), .A2(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n345), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n367), .A2(new_n332), .B1(new_n346), .B2(new_n349), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(KEYINPUT85), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n369), .A3(KEYINPUT4), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n363), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n331), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT82), .B1(new_n326), .B2(new_n331), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n346), .A2(new_n349), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n348), .A2(new_n347), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n365), .B2(new_n366), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n339), .A2(new_n350), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n370), .A2(new_n372), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n373), .A2(new_n374), .A3(new_n368), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n369), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  INV_X1    g191(.A(new_n314), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n361), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n323), .A2(new_n324), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n355), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n329), .A2(new_n313), .A3(new_n330), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n331), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n379), .A3(new_n399), .A4(new_n381), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n384), .ZN(new_n401));
  INV_X1    g200(.A(new_n371), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n351), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT84), .B1(new_n351), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n351), .A2(new_n352), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT85), .B1(new_n363), .B2(new_n368), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n401), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n387), .B1(new_n391), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(G57gat), .B(G85gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n387), .B(new_n415), .C1(new_n391), .C2(new_n410), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(KEYINPUT86), .A3(new_n418), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n417), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n419), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(KEYINPUT87), .A3(new_n424), .A4(new_n417), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n311), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT33), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n276), .A2(new_n363), .A3(new_n278), .A4(new_n279), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT68), .B1(new_n291), .B2(new_n229), .ZN(new_n436));
  INV_X1    g235(.A(new_n279), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(KEYINPUT72), .A3(new_n363), .A4(new_n276), .ZN(new_n439));
  INV_X1    g238(.A(new_n363), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n280), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT64), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n442), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n432), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G71gat), .B(G99gat), .Z(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n442), .A2(new_n445), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n431), .B1(new_n451), .B2(KEYINPUT33), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT74), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT74), .B(new_n457), .C1(new_n446), .C2(new_n447), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n452), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n442), .A2(KEYINPUT34), .A3(new_n445), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n435), .A2(new_n439), .A3(new_n441), .A4(new_n444), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n464), .A2(KEYINPUT75), .A3(KEYINPUT34), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT75), .B1(new_n464), .B2(KEYINPUT34), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n457), .B1(new_n446), .B2(new_n447), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  INV_X1    g271(.A(new_n467), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n452), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G50gat), .ZN(new_n475));
  INV_X1    g274(.A(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n380), .B1(new_n212), .B2(new_n286), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n376), .B2(new_n378), .ZN(new_n479));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n286), .B1(new_n368), .B2(new_n380), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n479), .B(new_n480), .C1(new_n294), .C2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n213), .B2(new_n217), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n215), .A2(new_n267), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n368), .B1(new_n484), .B2(new_n380), .ZN(new_n485));
  OAI211_X1 g284(.A(G228gat), .B(G233gat), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G22gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n482), .B2(new_n486), .ZN(new_n490));
  OAI21_X1  g289(.A(G78gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(G78gat), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(KEYINPUT88), .A3(new_n493), .A4(new_n488), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n477), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n494), .A3(new_n477), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n468), .A2(new_n474), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n430), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT35), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n306), .A2(new_n503), .A3(new_n310), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n468), .A2(new_n504), .A3(new_n474), .A4(new_n498), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI221_X4 g308(.A(new_n467), .B1(new_n448), .B2(new_n451), .C1(new_n471), .C2(new_n459), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n473), .B1(new_n472), .B2(new_n452), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT36), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n468), .A2(new_n513), .A3(new_n474), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n303), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n295), .B1(new_n300), .B2(new_n294), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT89), .B1(new_n519), .B2(KEYINPUT37), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n204), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n281), .A2(new_n218), .A3(new_n283), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n293), .B2(new_n294), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n501), .A2(new_n309), .A3(new_n502), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT38), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(KEYINPUT37), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n389), .A2(new_n388), .A3(new_n385), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(KEYINPUT39), .C1(new_n384), .C2(new_n383), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n383), .A2(KEYINPUT39), .A3(new_n384), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n415), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT40), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n417), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n537), .B2(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n311), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n498), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n532), .A2(new_n541), .B1(new_n429), .B2(new_n498), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n509), .B1(new_n515), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  AOI21_X1  g344(.A(G1gat), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n546), .B(new_n548), .Z(new_n549));
  XOR2_X1   g348(.A(KEYINPUT94), .B(G8gat), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n546), .B(new_n548), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G8gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G29gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n564));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n555), .A2(KEYINPUT96), .A3(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n555), .B2(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT13), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n568), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT95), .B1(new_n579), .B2(new_n555), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n568), .B(KEYINPUT17), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n551), .A4(new_n554), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n573), .A2(new_n580), .A3(new_n583), .A4(new_n575), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n577), .B(new_n590), .C1(new_n585), .C2(new_n584), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G169gat), .B(G197gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT92), .ZN(new_n594));
  XOR2_X1   g393(.A(G113gat), .B(G141gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT91), .B(KEYINPUT11), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT12), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n589), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n591), .B(new_n599), .C1(new_n586), .C2(new_n588), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n543), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G232gat), .ZN(new_n614));
  INV_X1    g413(.A(G233gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n568), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n579), .B2(new_n613), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(KEYINPUT99), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(KEYINPUT99), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n618), .B(new_n626), .C1(KEYINPUT99), .C2(new_n619), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n622), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n622), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(G64gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(G57gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G71gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n493), .ZN(new_n638));
  NOR2_X1   g437(.A1(G71gat), .A2(G78gat), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n638), .A2(new_n639), .B1(new_n632), .B2(KEYINPUT98), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n322), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n555), .B1(KEYINPUT21), .B2(new_n641), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G155gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n613), .B(new_n641), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n641), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n657), .B2(new_n656), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n661), .A2(KEYINPUT100), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n661), .B2(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n631), .A2(new_n654), .A3(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n427), .A2(new_n428), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n604), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  INV_X1    g479(.A(new_n311), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n672), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n543), .A2(new_n603), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n683), .A2(KEYINPUT103), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n683), .B2(G8gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n685), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI211_X1 g493(.A(KEYINPUT104), .B(new_n686), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(G1325gat));
  NAND2_X1  g495(.A1(new_n604), .A2(new_n673), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT36), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n513), .B1(new_n468), .B2(new_n474), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n512), .A2(KEYINPUT105), .A3(new_n514), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n510), .A2(new_n511), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n672), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n604), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(G1326gat));
  NOR2_X1   g508(.A1(new_n697), .A2(new_n498), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(new_n603), .ZN(new_n713));
  INV_X1    g512(.A(new_n668), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(new_n654), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n543), .A2(new_n630), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n560), .A3(new_n678), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n505), .A2(new_n506), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n705), .A2(KEYINPUT90), .A3(new_n498), .A4(new_n504), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n429), .A3(new_n498), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(KEYINPUT35), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n542), .A2(new_n515), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT44), .B(new_n630), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n715), .B(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n491), .A2(new_n494), .A3(new_n477), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n495), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n526), .B1(new_n521), .B2(new_n524), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n521), .A2(new_n530), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n529), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n539), .B2(new_n311), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n430), .A2(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n512), .A2(KEYINPUT105), .A3(new_n514), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT105), .B1(new_n512), .B2(new_n514), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n631), .B1(new_n737), .B2(new_n509), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n725), .B(new_n727), .C1(new_n738), .C2(KEYINPUT44), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n542), .B1(new_n701), .B2(new_n702), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n630), .B1(new_n742), .B2(new_n723), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n745), .A2(KEYINPUT107), .A3(new_n725), .A4(new_n727), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n741), .A2(new_n678), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n719), .B1(new_n560), .B2(new_n747), .ZN(G1328gat));
  NAND3_X1  g547(.A1(new_n741), .A2(new_n311), .A3(new_n746), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G36gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n681), .A2(G36gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n717), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n755));
  INV_X1    g554(.A(new_n753), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n716), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n750), .A2(KEYINPUT109), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1329gat));
  NOR3_X1   g562(.A1(new_n716), .A2(G43gat), .A3(new_n706), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G43gat), .B1(new_n739), .B2(new_n703), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n741), .A2(new_n702), .A3(new_n746), .A4(new_n701), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(G43gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g570(.A1(new_n716), .A2(G50gat), .A3(new_n498), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT48), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G50gat), .B1(new_n739), .B2(new_n498), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n741), .A2(new_n729), .A3(new_n746), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n772), .B1(new_n777), .B2(G50gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g578(.A(new_n654), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n630), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n713), .A2(new_n781), .A3(new_n714), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n737), .B2(new_n509), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n678), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g584(.A(new_n681), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT110), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1333gat));
  OR2_X1    g589(.A1(new_n705), .A2(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n705), .A2(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(G71gat), .B1(new_n783), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n703), .A2(new_n637), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g596(.A1(new_n783), .A2(new_n729), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n603), .A2(new_n654), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n714), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT112), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n745), .A2(new_n725), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n677), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(KEYINPUT113), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n804), .B2(KEYINPUT113), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n738), .A2(new_n807), .A3(new_n800), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n630), .B(new_n800), .C1(new_n742), .C2(new_n723), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n678), .A2(new_n608), .A3(new_n714), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n805), .A2(new_n806), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  OAI21_X1  g612(.A(G92gat), .B1(new_n803), .B2(new_n681), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n681), .A2(new_n668), .A3(G92gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n814), .B(new_n815), .C1(new_n811), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n809), .B2(KEYINPUT114), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n807), .B2(KEYINPUT115), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n820), .A2(new_n807), .B1(new_n809), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n816), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n814), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n825), .B2(new_n815), .ZN(G1337gat));
  OAI21_X1  g625(.A(G99gat), .B1(new_n803), .B2(new_n703), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n706), .A2(G99gat), .A3(new_n668), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n811), .B2(new_n828), .ZN(G1338gat));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n820), .A2(new_n807), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n809), .A2(new_n822), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n498), .A2(new_n668), .A3(G106gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n745), .A2(new_n729), .A3(new_n725), .A4(new_n802), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n808), .A2(new_n810), .A3(new_n834), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n830), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n831), .A3(new_n839), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n823), .A2(new_n834), .B1(G106gat), .B2(new_n836), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT116), .B(new_n842), .C1(new_n843), .C2(new_n831), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n327), .A2(new_n328), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n669), .A2(new_n603), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n658), .A2(new_n659), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n655), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n658), .A2(new_n659), .A3(new_n656), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n664), .B1(new_n660), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT117), .A4(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n661), .A2(new_n664), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n854), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n857), .A2(new_n630), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n573), .A2(new_n583), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n575), .B1(new_n864), .B2(new_n580), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n574), .A2(new_n576), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n598), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(KEYINPUT18), .A3(new_n575), .A4(new_n580), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n577), .A3(new_n587), .A4(new_n600), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n848), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AND4_X1   g670(.A1(new_n860), .A2(new_n862), .A3(new_n856), .A4(new_n855), .ZN(new_n872));
  INV_X1    g671(.A(new_n870), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(KEYINPUT118), .A3(new_n630), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n870), .A2(new_n668), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n603), .B2(new_n872), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n871), .B(new_n874), .C1(new_n876), .C2(new_n630), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n847), .B1(new_n877), .B2(new_n780), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n499), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n677), .A2(new_n311), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n603), .ZN(new_n882));
  MUX2_X1   g681(.A(new_n846), .B(G113gat), .S(new_n882), .Z(G1340gat));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n714), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n654), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n354), .A2(new_n316), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1342gat));
  NAND2_X1  g687(.A1(new_n880), .A2(new_n630), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n891), .B(new_n892), .Z(G1343gat));
  NAND2_X1  g692(.A1(new_n860), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n858), .A2(new_n895), .A3(new_n859), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n857), .A2(new_n894), .A3(new_n862), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n601), .B2(new_n602), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n631), .B1(new_n898), .B2(new_n875), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n874), .A2(new_n871), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n847), .B1(new_n901), .B2(new_n780), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n498), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n877), .A2(new_n780), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n904), .B(new_n729), .C1(new_n905), .C2(new_n847), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n703), .A2(new_n880), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n603), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G141gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n878), .A2(new_n498), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n603), .A2(new_n343), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n340), .A3(new_n714), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n668), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .A3(new_n340), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT57), .B1(new_n878), .B2(new_n498), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n498), .A2(KEYINPUT57), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n872), .A2(new_n630), .A3(new_n873), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n654), .B1(new_n899), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n672), .A2(new_n603), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n714), .A3(new_n907), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n921), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n917), .B1(new_n920), .B2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n918), .B2(new_n780), .ZN(new_n932));
  INV_X1    g731(.A(G155gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n933), .A3(new_n654), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1346gat));
  NOR2_X1   g734(.A1(new_n889), .A2(G162gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n910), .A2(new_n703), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  OAI21_X1  g737(.A(G162gat), .B1(new_n918), .B2(new_n631), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n678), .A2(new_n681), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n879), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n221), .A3(new_n603), .ZN(new_n944));
  INV_X1    g743(.A(new_n878), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n729), .B1(new_n791), .B2(new_n792), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(new_n713), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(G169gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n948), .B2(G169gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n944), .B1(new_n950), .B2(new_n951), .ZN(G1348gat));
  OAI21_X1  g751(.A(G176gat), .B1(new_n947), .B2(new_n668), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n714), .A2(new_n222), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n942), .B2(new_n954), .ZN(G1349gat));
  NAND2_X1  g754(.A1(new_n238), .A2(G183gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n654), .A2(new_n956), .A3(new_n288), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n943), .A2(KEYINPUT123), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n942), .B2(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n963), .A2(KEYINPUT60), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n654), .A3(new_n941), .A4(new_n946), .ZN(new_n965));
  INV_X1    g764(.A(new_n261), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n965), .A2(new_n966), .B1(new_n963), .B2(KEYINPUT60), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n962), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n962), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n943), .A2(new_n233), .A3(new_n630), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n947), .A2(new_n631), .ZN(new_n972));
  XNOR2_X1  g771(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(G190gat), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n972), .B2(G190gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  NAND3_X1  g775(.A1(new_n703), .A2(new_n311), .A3(new_n729), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n878), .A2(new_n678), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n603), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n941), .A2(new_n703), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n928), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n713), .A2(new_n205), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n982), .A2(new_n206), .A3(new_n714), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n928), .A2(new_n714), .A3(new_n984), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n989), .B(new_n990), .C1(new_n206), .C2(new_n991), .ZN(G1353gat));
  OR3_X1    g791(.A1(new_n981), .A2(G211gat), .A3(new_n780), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n922), .A2(new_n927), .A3(new_n654), .A4(new_n984), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT127), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1354gat));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n630), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G218gat), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n631), .A2(G218gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n981), .B2(new_n1004), .ZN(G1355gat));
endmodule


