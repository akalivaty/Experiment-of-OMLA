//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  XOR2_X1   g0004(.A(KEYINPUT65), .B(G77), .Z(new_n205));
  INV_X1    g0005(.A(G244), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n204), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n204), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n214), .B(new_n217), .C1(new_n220), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  INV_X1    g0041(.A(G13), .ZN(new_n242));
  NOR3_X1   g0042(.A1(new_n242), .A2(new_n219), .A3(G1), .ZN(new_n243));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n218), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(G50), .B1(new_n219), .B2(G1), .ZN(new_n248));
  INV_X1    g0048(.A(new_n243), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n247), .A2(new_n248), .B1(G50), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(KEYINPUT8), .B(G58), .Z(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n219), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G50), .A2(G58), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n219), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OR3_X1    g0061(.A1(new_n254), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n250), .B1(new_n262), .B2(new_n245), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n265));
  INV_X1    g0065(.A(G190), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n273), .B(new_n274), .C1(new_n205), .C2(new_n271), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G274), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n276), .B2(new_n278), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT66), .A3(new_n285), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n285), .B1(new_n276), .B2(new_n278), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G226), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n282), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(G200), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n296), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  AOI211_X1 g0104(.A(new_n263), .B(new_n303), .C1(new_n304), .C2(new_n296), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G232), .A2(G1698), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n272), .A2(G238), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n271), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n281), .B(new_n308), .C1(G107), .C2(new_n271), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n294), .A2(G244), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n293), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(new_n266), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(G200), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n253), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n252), .A2(new_n259), .B1(new_n219), .B2(new_n205), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n245), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  INV_X1    g0119(.A(G1), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n246), .A2(new_n321), .B1(new_n205), .B2(new_n243), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n312), .A2(new_n313), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n311), .A2(G179), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n311), .A2(new_n304), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n302), .A2(new_n305), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n293), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n292), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n227), .A2(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G226), .B2(G1698), .ZN(new_n334));
  AND2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G97), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n334), .A2(new_n337), .B1(new_n268), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n281), .B1(G238), .B2(new_n294), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n331), .A2(KEYINPUT13), .A3(new_n340), .A4(new_n332), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(G200), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n346), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n331), .A2(new_n332), .A3(new_n340), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n266), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT72), .B1(new_n249), .B2(G68), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n351), .B(KEYINPUT12), .Z(new_n352));
  OAI211_X1 g0152(.A(new_n246), .B(G68), .C1(G1), .C2(new_n219), .ZN(new_n353));
  INV_X1    g0153(.A(G50), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n259), .A2(new_n354), .B1(new_n219), .B2(G68), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n253), .A2(new_n319), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n245), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT11), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n345), .A2(new_n350), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n343), .A2(G169), .A3(new_n344), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n343), .A2(new_n363), .A3(G169), .A4(new_n344), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n349), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n360), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n271), .B2(G20), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n256), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G58), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n256), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n221), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n259), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n369), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT74), .B(new_n369), .C1(new_n373), .C2(new_n378), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n271), .A2(new_n370), .A3(G20), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n337), .B2(new_n219), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n376), .B(KEYINPUT73), .C1(new_n377), .C2(new_n259), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT16), .A4(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n381), .A2(new_n245), .A3(new_n382), .A4(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n252), .B1(new_n320), .B2(G20), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n246), .B1(new_n243), .B2(new_n252), .ZN(new_n392));
  OR2_X1    g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G226), .B2(new_n272), .ZN(new_n394));
  INV_X1    g0194(.A(G87), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n394), .A2(new_n337), .B1(new_n268), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n281), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n294), .A2(G232), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(G190), .A3(new_n293), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n293), .A3(new_n398), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G200), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n390), .A2(new_n392), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n390), .A2(new_n392), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(G179), .A3(new_n293), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(G169), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n329), .A2(new_n368), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n243), .A2(new_n338), .ZN(new_n417));
  INV_X1    g0217(.A(new_n245), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n320), .A2(G33), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n249), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n338), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n371), .A2(new_n372), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(G107), .B1(G77), .B2(new_n258), .ZN(new_n424));
  NOR2_X1   g0224(.A1(G97), .A2(G107), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT6), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(KEYINPUT6), .B2(new_n338), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT75), .B(G107), .Z(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  OAI21_X1  g0230(.A(G20), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n418), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(KEYINPUT4), .A2(G244), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n272), .B(new_n433), .C1(new_n335), .C2(new_n336), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G283), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n206), .B1(new_n269), .B2(new_n270), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n434), .B(new_n435), .C1(new_n436), .C2(KEYINPUT4), .ZN(new_n437));
  OAI21_X1  g0237(.A(G250), .B1(new_n335), .B2(new_n336), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n272), .B1(new_n438), .B2(KEYINPUT4), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n281), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n283), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT76), .B1(new_n283), .B2(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G41), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n283), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(KEYINPUT77), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n284), .A2(G1), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(G41), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n444), .A2(new_n291), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n448), .A3(new_n450), .A4(new_n451), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(G257), .A3(new_n286), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n440), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n422), .B(new_n432), .C1(G200), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT79), .ZN(new_n458));
  AND4_X1   g0258(.A1(KEYINPUT78), .A2(new_n440), .A3(new_n453), .A4(new_n455), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n453), .A2(new_n455), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT78), .B1(new_n460), .B2(new_n440), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n462), .B2(G190), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT79), .A4(new_n266), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n432), .A2(new_n422), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n456), .A2(G179), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n304), .B1(new_n459), .B2(new_n461), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n447), .A2(new_n448), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n450), .A2(new_n451), .ZN(new_n473));
  OAI211_X1 g0273(.A(G270), .B(new_n286), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n454), .A2(KEYINPUT82), .A3(G270), .A4(new_n286), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G264), .B(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(new_n272), .C1(new_n335), .C2(new_n336), .ZN(new_n480));
  INV_X1    g0280(.A(G303), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n271), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n281), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n453), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n435), .B(new_n219), .C1(G33), .C2(new_n338), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n245), .C1(new_n219), .C2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n249), .A2(G116), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n420), .B2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(G169), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G179), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n482), .B2(new_n281), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n478), .A2(new_n453), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n492), .A2(new_n493), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n491), .B1(new_n484), .B2(G200), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n266), .B2(new_n484), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT25), .B1(new_n243), .B2(new_n503), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n421), .A2(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n219), .B(G87), .C1(new_n335), .C2(new_n336), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n271), .A2(new_n510), .A3(new_n219), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(KEYINPUT23), .C1(new_n219), .C2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n503), .A2(G20), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(KEYINPUT23), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n503), .A3(G20), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n512), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n245), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT84), .B(new_n245), .C1(new_n524), .C2(new_n525), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n507), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n454), .A2(G264), .A3(new_n286), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT85), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n454), .A2(new_n533), .A3(G264), .A4(new_n286), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n271), .A2(G250), .A3(new_n272), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G294), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n532), .A2(new_n534), .B1(new_n538), .B2(new_n281), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n453), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n304), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G179), .B2(new_n540), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  INV_X1    g0344(.A(G200), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n540), .A2(G190), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n540), .A2(new_n544), .A3(G190), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n530), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G250), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n284), .B2(G1), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n320), .A2(new_n290), .A3(G45), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n286), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n556));
  OAI211_X1 g0356(.A(G238), .B(new_n272), .C1(new_n335), .C2(new_n336), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n559), .B2(new_n281), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(KEYINPUT80), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT80), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n562), .B(new_n555), .C1(new_n559), .C2(new_n281), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n271), .A2(new_n219), .A3(G68), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n253), .A2(new_n338), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(KEYINPUT19), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g0368(.A(KEYINPUT81), .B(G87), .Z(new_n569));
  NAND3_X1  g0369(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(new_n425), .B1(new_n219), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n245), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n315), .A2(new_n243), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(G87), .B2(new_n420), .ZN(new_n575));
  OAI21_X1  g0375(.A(G200), .B1(new_n561), .B2(new_n563), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n565), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n564), .A2(new_n495), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n304), .B1(new_n561), .B2(new_n563), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n572), .B(new_n573), .C1(new_n315), .C2(new_n421), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n502), .A2(new_n543), .A3(new_n550), .A4(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n416), .A2(new_n471), .A3(new_n583), .ZN(G372));
  INV_X1    g0384(.A(new_n302), .ZN(new_n585));
  INV_X1    g0385(.A(new_n360), .ZN(new_n586));
  INV_X1    g0386(.A(new_n327), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n367), .B2(new_n359), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n411), .B(new_n413), .C1(new_n588), .C2(new_n405), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n305), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT26), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n582), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n560), .A2(new_n545), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT87), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n565), .A3(new_n575), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n494), .B(new_n499), .C1(new_n530), .C2(new_n542), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n465), .A2(new_n598), .A3(new_n550), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(new_n470), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n593), .B1(new_n600), .B2(KEYINPUT26), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n578), .B(new_n580), .C1(G169), .C2(new_n560), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n590), .B1(new_n416), .B2(new_n604), .ZN(G369));
  AND2_X1   g0405(.A1(new_n543), .A2(new_n550), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n320), .A2(new_n219), .A3(G13), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(KEYINPUT27), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT88), .ZN(new_n609));
  INV_X1    g0409(.A(G213), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n607), .B2(KEYINPUT27), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(G343), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT89), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT89), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n606), .B1(new_n530), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n543), .B2(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n491), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n502), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n494), .A2(new_n499), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G330), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n543), .A2(new_n615), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n621), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(G399));
  INV_X1    g0429(.A(new_n215), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(G41), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n224), .ZN(new_n632));
  INV_X1    g0432(.A(G116), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n569), .A2(new_n633), .A3(new_n425), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G1), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT28), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n560), .A2(G179), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n540), .A2(new_n638), .A3(new_n456), .A4(new_n484), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n497), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT77), .B1(new_n447), .B2(new_n448), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n286), .A2(G274), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n643), .A2(new_n644), .A3(new_n473), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n476), .A2(new_n477), .B1(new_n449), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(KEYINPUT90), .A3(new_n496), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n532), .A2(new_n534), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n538), .A2(new_n281), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(new_n561), .A3(new_n563), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n648), .A2(new_n462), .A3(KEYINPUT30), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT92), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT78), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n456), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n460), .A2(KEYINPUT78), .A3(new_n440), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n656), .A2(new_n564), .A3(new_n657), .A4(new_n539), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT30), .A4(new_n648), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n640), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n648), .A2(new_n462), .A3(new_n652), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT30), .B1(new_n662), .B2(KEYINPUT91), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n648), .A2(new_n462), .A3(new_n664), .A4(new_n652), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT93), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n497), .A2(new_n641), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT90), .B1(new_n646), .B2(new_n496), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n656), .A2(new_n564), .A3(new_n657), .A4(new_n539), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT91), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  AND4_X1   g0472(.A1(KEYINPUT93), .A2(new_n671), .A3(new_n672), .A4(new_n665), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n661), .B1(new_n666), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT31), .B1(new_n674), .B2(new_n615), .ZN(new_n675));
  INV_X1    g0475(.A(new_n471), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n577), .A2(new_n581), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(new_n606), .A3(new_n679), .A4(new_n616), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n663), .A2(new_n665), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n661), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n616), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(G330), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n615), .B1(new_n601), .B2(new_n602), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n602), .A2(new_n596), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT94), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n592), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT94), .B1(new_n691), .B2(new_n591), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n678), .B2(new_n470), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n602), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n692), .A2(new_n465), .A3(new_n470), .A4(new_n550), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n616), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n688), .B1(new_n690), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n637), .B1(new_n707), .B2(G1), .ZN(G364));
  NOR2_X1   g0508(.A1(new_n242), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n320), .B1(new_n709), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n631), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n624), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G330), .B2(new_n622), .ZN(new_n714));
  INV_X1    g0514(.A(new_n712), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n218), .B1(G20), .B2(new_n304), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT97), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n266), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G326), .ZN(new_n722));
  NAND2_X1  g0522(.A1(G20), .A2(G179), .ZN(new_n723));
  AOI21_X1  g0523(.A(G200), .B1(new_n723), .B2(KEYINPUT96), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(KEYINPUT96), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G311), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n721), .A2(new_n722), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n719), .A2(G190), .ZN(new_n730));
  XNOR2_X1  g0530(.A(KEYINPUT33), .B(G317), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n545), .A2(G179), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G20), .A3(G190), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n337), .B1(new_n734), .B2(new_n481), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n219), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G329), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n737), .A2(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n735), .B(new_n742), .C1(G294), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n725), .A2(new_n266), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n732), .B(new_n745), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n205), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n720), .A2(G50), .B1(new_n726), .B2(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n730), .A2(G68), .B1(new_n747), .B2(G58), .ZN(new_n752));
  INV_X1    g0552(.A(new_n744), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n338), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n569), .A2(new_n734), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n271), .B1(new_n737), .B2(new_n503), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n740), .A2(new_n377), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n751), .A2(new_n752), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n717), .B1(new_n749), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n215), .A2(G355), .A3(new_n271), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n630), .A2(new_n271), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n223), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n237), .A2(G45), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n766), .B1(G116), .B2(new_n215), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n715), .B(new_n761), .C1(new_n765), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n764), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n622), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n714), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  NAND2_X1  g0575(.A1(new_n615), .A2(new_n325), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n587), .B1(new_n776), .B2(new_n323), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n327), .A2(new_n615), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n689), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n712), .B1(new_n780), .B2(new_n687), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n687), .B2(new_n780), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G137), .A2(new_n720), .B1(new_n730), .B2(G150), .ZN(new_n783));
  INV_X1    g0583(.A(G143), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n784), .B2(new_n748), .C1(new_n377), .C2(new_n727), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  NOR2_X1   g0586(.A1(new_n753), .A2(new_n374), .ZN(new_n787));
  INV_X1    g0587(.A(G132), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n271), .B1(new_n740), .B2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n734), .A2(new_n354), .B1(new_n737), .B2(new_n256), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n786), .A2(new_n787), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n740), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n271), .B1(new_n792), .B2(G311), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n395), .B2(new_n737), .C1(new_n503), .C2(new_n734), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n754), .B(new_n794), .C1(G303), .C2(new_n720), .ZN(new_n795));
  INV_X1    g0595(.A(new_n730), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n796), .A2(new_n738), .B1(new_n727), .B2(new_n633), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(KEYINPUT98), .B2(new_n797), .C1(new_n798), .C2(new_n748), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(KEYINPUT98), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n716), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n716), .A2(new_n762), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n715), .B1(new_n319), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(new_n763), .C2(new_n779), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  NOR2_X1   g0606(.A1(new_n709), .A2(new_n320), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT40), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n369), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(new_n245), .A3(new_n389), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT101), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n811), .A2(new_n812), .A3(new_n392), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n811), .B2(new_n392), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n609), .A2(new_n611), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n409), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n403), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT37), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n406), .A2(new_n816), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n410), .A2(new_n821), .A3(new_n822), .A4(new_n403), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n405), .B2(new_n414), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n826), .A3(KEYINPUT38), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT38), .B1(new_n824), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n615), .A2(new_n359), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n368), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n360), .B2(new_n367), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(KEYINPUT100), .B(new_n834), .C1(new_n360), .C2(new_n367), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n833), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n779), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n654), .A2(new_n660), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n639), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT93), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n681), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n663), .A2(KEYINPUT93), .A3(new_n665), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n683), .B1(new_n846), .B2(new_n616), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n583), .A2(new_n471), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n674), .A2(new_n684), .B1(new_n848), .B2(new_n616), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n840), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n831), .B1(new_n850), .B2(KEYINPUT102), .ZN(new_n851));
  INV_X1    g0651(.A(new_n779), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n368), .A2(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n838), .ZN(new_n854));
  INV_X1    g0654(.A(new_n684), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n680), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n856), .B2(new_n675), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n808), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT103), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n406), .B(new_n816), .C1(new_n405), .C2(new_n414), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n410), .A2(new_n821), .A3(new_n403), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n823), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n808), .B1(new_n869), .B2(new_n827), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n850), .B2(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n860), .B1(new_n862), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n416), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n847), .A2(new_n849), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(G330), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n839), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n603), .A2(new_n616), .A3(new_n779), .ZN(new_n880));
  INV_X1    g0680(.A(new_n778), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n831), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT39), .B1(new_n869), .B2(new_n827), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(KEYINPUT39), .B2(new_n830), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n367), .A2(new_n359), .A3(new_n616), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n414), .A2(new_n815), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n690), .A2(new_n706), .A3(new_n873), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n590), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n807), .B1(new_n878), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n878), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n220), .A2(G116), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n429), .A2(new_n430), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(KEYINPUT35), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(KEYINPUT35), .B2(new_n898), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n223), .A2(new_n375), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n902), .A2(new_n205), .B1(G50), .B2(new_n256), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n242), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT99), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n895), .A2(new_n906), .ZN(G367));
  INV_X1    g0707(.A(new_n767), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n765), .B1(new_n215), .B2(new_n315), .C1(new_n908), .C2(new_n233), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n712), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n616), .A2(new_n575), .ZN(new_n911));
  INV_X1    g0711(.A(new_n602), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n691), .B2(new_n911), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n721), .A2(new_n784), .B1(new_n748), .B2(new_n260), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G50), .B2(new_n726), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n730), .A2(G159), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n753), .A2(new_n256), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(KEYINPUT109), .B(G137), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n734), .A2(new_n374), .B1(new_n740), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n737), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n337), .B(new_n921), .C1(new_n750), .C2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n916), .A2(new_n917), .A3(new_n919), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n734), .A2(new_n633), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT46), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n730), .A2(G294), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n337), .B1(new_n737), .B2(new_n338), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(G317), .B2(new_n792), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n720), .A2(G311), .B1(new_n747), .B2(G303), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n927), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n726), .A2(G283), .B1(G107), .B2(new_n744), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT108), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n924), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  OAI221_X1 g0735(.A(new_n910), .B1(new_n914), .B2(new_n772), .C1(new_n935), .C2(new_n717), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n914), .B(KEYINPUT43), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n470), .A2(new_n616), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT104), .Z(new_n940));
  OAI21_X1  g0740(.A(new_n676), .B1(new_n466), .B2(new_n616), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n628), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT42), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT105), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n470), .B1(new_n942), .B2(new_n543), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n616), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n938), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n950), .B2(KEYINPUT106), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n952), .A2(new_n955), .B1(new_n625), .B2(new_n942), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n625), .A2(new_n942), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(new_n951), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n628), .A2(new_n626), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n942), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT44), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n942), .A2(new_n961), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n624), .A3(new_n618), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n625), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n628), .B1(new_n618), .B2(new_n627), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n624), .A2(KEYINPUT107), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n623), .B(KEYINPUT107), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n707), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n707), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n631), .B(KEYINPUT41), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n711), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n936), .B1(new_n960), .B2(new_n978), .ZN(G387));
  OR2_X1    g0779(.A1(new_n618), .A2(new_n772), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n230), .A2(new_n284), .A3(new_n271), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n284), .B1(new_n256), .B2(new_n319), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n252), .B2(G50), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n251), .A2(KEYINPUT50), .A3(new_n354), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n634), .B1(new_n986), .B2(new_n271), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n630), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n765), .B1(new_n215), .B2(new_n503), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n712), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n721), .A2(new_n377), .B1(new_n748), .B2(new_n354), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G68), .B2(new_n726), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n730), .A2(new_n251), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n315), .A2(new_n753), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n271), .B1(new_n737), .B2(new_n338), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n205), .A2(new_n734), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(G150), .C2(new_n792), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n753), .A2(new_n738), .B1(new_n734), .B2(new_n798), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G303), .A2(new_n726), .B1(new_n747), .B2(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n728), .B2(new_n796), .C1(new_n746), .C2(new_n721), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT49), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n337), .B1(new_n740), .B2(new_n722), .C1(new_n633), .C2(new_n737), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT110), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n990), .B1(new_n1008), .B2(new_n716), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n974), .A2(new_n711), .B1(new_n980), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n707), .A2(new_n974), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n631), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n707), .B2(new_n974), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1013), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(G393));
  NOR2_X1   g0818(.A1(new_n908), .A2(new_n240), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n765), .B1(new_n215), .B2(new_n338), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n712), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n720), .A2(G317), .B1(new_n747), .B2(G311), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n337), .B1(new_n737), .B2(new_n503), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n734), .A2(new_n738), .B1(new_n740), .B2(new_n746), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G116), .C2(new_n744), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n798), .B2(new_n727), .C1(new_n481), .C2(new_n796), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n271), .B1(new_n737), .B2(new_n395), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n734), .A2(new_n256), .B1(new_n740), .B2(new_n784), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G77), .C2(new_n744), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n354), .B2(new_n796), .C1(new_n252), .C2(new_n727), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n720), .A2(G150), .B1(new_n747), .B2(G159), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT51), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1023), .A2(new_n1027), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1021), .B1(new_n1034), .B2(new_n716), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n942), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n772), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n967), .A3(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(new_n975), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n631), .B1(new_n969), .B2(new_n975), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1037), .B1(new_n710), .B2(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(G390));
  INV_X1    g0843(.A(G330), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n847), .B2(new_n849), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n879), .B1(new_n1046), .B2(new_n852), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n881), .B1(new_n704), .B2(new_n777), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n779), .C1(new_n675), .C2(new_n686), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(new_n879), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1047), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n854), .A2(new_n1045), .B1(new_n1050), .B2(new_n879), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n778), .B1(new_n689), .B2(new_n779), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(KEYINPUT114), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT114), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1050), .A2(new_n879), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n854), .B(G330), .C1(new_n856), .C2(new_n675), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1055), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1053), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1046), .A2(new_n416), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n892), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1059), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n615), .B(new_n852), .C1(new_n601), .C2(new_n602), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n839), .B1(new_n1068), .B2(new_n778), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n885), .B1(new_n1069), .B2(new_n886), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT38), .B1(new_n863), .B2(new_n866), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n886), .B1(new_n828), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1048), .B2(new_n839), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1067), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n869), .A2(new_n827), .ZN(new_n1075));
  MUX2_X1   g0875(.A(new_n1075), .B(new_n830), .S(KEYINPUT39), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n882), .B2(new_n887), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1073), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n1052), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1066), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n886), .B1(new_n1055), .B2(new_n879), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1051), .B(new_n1073), .C1(new_n1084), .C2(new_n1076), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1059), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n891), .B(new_n590), .C1(new_n416), .C2(new_n1046), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT114), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1060), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1091), .B2(new_n1053), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1014), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1087), .A2(new_n711), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1076), .A2(new_n762), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n734), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(G87), .B1(new_n792), .B2(G294), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n271), .B1(new_n922), .B2(G68), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n319), .B2(new_n753), .C1(new_n633), .C2(new_n748), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n730), .A2(G107), .B1(new_n726), .B2(G97), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n738), .B2(new_n721), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  AOI22_X1  g0904(.A1(new_n720), .A2(G128), .B1(new_n726), .B2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n788), .B2(new_n748), .C1(new_n796), .C2(new_n920), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n734), .A2(new_n260), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n744), .A2(G159), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n922), .A2(G50), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n337), .B1(new_n792), .B2(G125), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1101), .A2(new_n1103), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n716), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n802), .A2(new_n252), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1096), .A2(new_n712), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1094), .A2(new_n1095), .A3(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1063), .A2(new_n1074), .A3(new_n1079), .A4(new_n1065), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n1065), .ZN(new_n1120));
  OAI21_X1  g0920(.A(G330), .B1(new_n871), .B2(new_n862), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n830), .B1(new_n857), .B2(new_n858), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT40), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT117), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT40), .B1(new_n828), .B2(new_n1071), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n857), .B2(new_n861), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1044), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n860), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n302), .A2(new_n305), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n263), .A2(new_n815), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT116), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1132), .B(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1125), .A2(new_n1131), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n1130), .A3(new_n860), .A4(new_n1129), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n890), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n890), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1139), .A2(new_n1143), .A3(new_n1140), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1120), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1120), .A2(new_n1142), .A3(KEYINPUT118), .A4(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1144), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1088), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1143), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT119), .B1(new_n1153), .B2(KEYINPUT57), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1118), .C1(new_n1156), .C2(new_n1151), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1149), .A2(new_n1154), .A3(new_n631), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n802), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n260), .B2(new_n753), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n730), .A2(G132), .B1(new_n726), .B2(G137), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n748), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(G125), .C2(new_n720), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n922), .A2(G159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n796), .A2(new_n338), .B1(new_n748), .B2(new_n503), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n737), .A2(new_n374), .B1(new_n740), .B2(new_n738), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n337), .A2(new_n283), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1173), .A2(new_n996), .A3(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n919), .C1(new_n315), .C2(new_n727), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1172), .B(new_n1176), .C1(G116), .C2(new_n720), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1174), .B(new_n354), .C1(G33), .C2(G41), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1180));
  AND4_X1   g0980(.A1(new_n1171), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n712), .B1(G50), .B2(new_n1159), .C1(new_n1181), .C2(new_n717), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1137), .B2(new_n762), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n711), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1158), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  NAND3_X1  g0987(.A1(new_n1091), .A2(new_n1088), .A3(new_n1053), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1066), .A2(new_n977), .A3(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT120), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n879), .A2(new_n762), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n712), .B1(G68), .B2(new_n1159), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n721), .A2(new_n788), .B1(new_n727), .B2(new_n260), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n730), .B2(new_n1104), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n271), .B1(new_n737), .B2(new_n374), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n734), .A2(new_n377), .B1(new_n740), .B2(new_n1163), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G50), .C2(new_n744), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1194), .B(new_n1197), .C1(new_n748), .C2(new_n920), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n734), .A2(new_n338), .B1(new_n740), .B2(new_n481), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  AOI22_X1  g1000(.A1(new_n720), .A2(G294), .B1(new_n747), .B2(G283), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n633), .C2(new_n796), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n271), .B1(new_n922), .B2(G77), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n994), .B(new_n1203), .C1(new_n503), .C2(new_n727), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1192), .B1(new_n1205), .B2(new_n716), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1063), .A2(new_n711), .B1(new_n1191), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1190), .A2(new_n1207), .ZN(G381));
  OR2_X1    g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(G384), .ZN(new_n1210));
  OR2_X1    g1010(.A1(G390), .A2(G387), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1210), .A2(new_n1211), .A3(G378), .A4(G381), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1186), .ZN(G407));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n610), .A2(G343), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1186), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(G213), .A3(new_n1216), .ZN(G409));
  NAND2_X1  g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(G390), .A2(G387), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT123), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(G390), .B2(G387), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1209), .B(new_n1218), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1209), .A2(new_n1218), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1211), .A2(new_n1224), .A3(new_n1221), .A4(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1158), .A2(G378), .A3(new_n1185), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1153), .A2(new_n977), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1185), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1214), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1215), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1188), .B(KEYINPUT60), .Z(new_n1232));
  NAND2_X1  g1032(.A1(new_n1066), .A2(new_n631), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1207), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(G384), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT62), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1215), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT125), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT125), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1240), .B(new_n1215), .C1(new_n1227), .C2(new_n1230), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1236), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1215), .A2(G2897), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1235), .B(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1226), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1242), .A2(KEYINPUT63), .A3(new_n1235), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT63), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1247), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1223), .A2(new_n1257), .A3(new_n1225), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1258), .A2(KEYINPUT124), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(KEYINPUT124), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1252), .A2(new_n1254), .A3(new_n1256), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1251), .A2(new_n1262), .ZN(G405));
  NAND2_X1  g1063(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1186), .A2(G378), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(new_n1235), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1235), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1226), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1226), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1264), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1226), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1264), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(G402));
endmodule


