//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n646, new_n649, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT66), .Z(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n470), .A2(G137), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n472), .B(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n470), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n479), .B1(new_n482), .B2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(G2105), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(KEYINPUT68), .A3(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT68), .B1(new_n484), .B2(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT69), .ZN(G162));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n472), .A2(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n470), .A3(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n499), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n472), .A3(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(G88), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G50), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(G75), .A2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n517), .B2(G62), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n513), .A2(KEYINPUT71), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n521), .A2(new_n522), .A3(new_n508), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n505), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n518), .A2(new_n519), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n521), .B2(new_n508), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT72), .A4(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n515), .A2(new_n532), .A3(new_n516), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n531), .A2(G63), .A3(G651), .A4(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n509), .A2(new_n510), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT6), .B(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n539), .A2(new_n542), .A3(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT75), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n538), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G168));
  INV_X1    g124(.A(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n540), .B2(new_n541), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G52), .A3(new_n539), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n536), .A2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(KEYINPUT76), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n531), .A2(G64), .A3(new_n533), .ZN(new_n558));
  INV_X1    g133(.A(G77), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n550), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n556), .A2(new_n557), .B1(G651), .B2(new_n560), .ZN(G171));
  NAND2_X1  g136(.A1(new_n551), .A2(new_n539), .ZN(new_n562));
  INV_X1    g137(.A(G43), .ZN(new_n563));
  INV_X1    g138(.A(new_n536), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT77), .B(G81), .Z(new_n565));
  OAI22_X1  g140(.A1(new_n562), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n531), .A2(G56), .A3(new_n533), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n519), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n535), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n536), .A2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n551), .A2(G53), .A3(new_n539), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n551), .A2(new_n584), .A3(G53), .A4(new_n539), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  NAND2_X1  g162(.A1(new_n560), .A2(G651), .ZN(new_n588));
  INV_X1    g163(.A(new_n557), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT76), .B1(new_n552), .B2(new_n553), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G301));
  NOR2_X1   g166(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT7), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n534), .B(new_n537), .C1(new_n592), .C2(new_n596), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n551), .A2(G51), .A3(new_n539), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT78), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n538), .A2(new_n544), .A3(new_n547), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G286));
  AND2_X1   g178(.A1(new_n531), .A2(new_n533), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n604), .B2(G74), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n543), .A2(G49), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n536), .A2(G87), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G288));
  NAND2_X1  g183(.A1(G48), .A2(G543), .ZN(new_n609));
  OR3_X1    g184(.A1(new_n508), .A2(KEYINPUT79), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT79), .B1(new_n508), .B2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n517), .A2(G61), .ZN(new_n613));
  AND2_X1   g188(.A1(G73), .A2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n536), .A2(G86), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(G305));
  NAND2_X1  g192(.A1(new_n536), .A2(G85), .ZN(new_n618));
  INV_X1    g193(.A(G47), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n562), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n531), .A2(G60), .A3(new_n533), .ZN(new_n621));
  NAND2_X1  g196(.A1(G72), .A2(G543), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n519), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n620), .B1(new_n624), .B2(KEYINPUT80), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n627), .ZN(G290));
  NAND2_X1  g203(.A1(G301), .A2(G868), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n517), .A2(new_n540), .A3(G92), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n551), .A2(G54), .A3(new_n539), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n633));
  INV_X1    g208(.A(G66), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n515), .B2(new_n516), .ZN(new_n635));
  AND2_X1   g210(.A1(G79), .A2(G543), .ZN(new_n636));
  OAI21_X1  g211(.A(G651), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n633), .B1(new_n632), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n631), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n629), .B1(new_n643), .B2(G868), .ZN(G284));
  OAI21_X1  g219(.A(new_n629), .B1(new_n643), .B2(G868), .ZN(G321));
  NOR2_X1   g220(.A1(G299), .A2(G868), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(G868), .B2(new_n602), .ZN(G297));
  AOI21_X1  g222(.A(new_n646), .B1(G868), .B2(new_n602), .ZN(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G868), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g228(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g229(.A1(new_n470), .A2(G2104), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n472), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n484), .A2(G135), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n482), .A2(G123), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n663), .A2(new_n470), .A3(G111), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n470), .B2(G111), .ZN(new_n665));
  OR2_X1    g240(.A1(G99), .A2(G2105), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G2104), .A3(new_n666), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n661), .B(new_n662), .C1(new_n664), .C2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2096), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(G2096), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n660), .A2(new_n669), .A3(new_n670), .ZN(G156));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2427), .B(G2430), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT14), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n673), .B2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1341), .B(G1348), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2451), .B(G2454), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT16), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(G14), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n687), .A2(KEYINPUT87), .A3(G14), .A4(new_n688), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G401));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  XOR2_X1   g270(.A(G2072), .B(G2078), .Z(new_n696));
  XOR2_X1   g271(.A(G2084), .B(G2090), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT18), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n696), .B(KEYINPUT17), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n698), .C1(new_n695), .C2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n695), .A3(new_n697), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G2096), .B(G2100), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G227));
  XOR2_X1   g282(.A(G1971), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT19), .ZN(new_n709));
  XOR2_X1   g284(.A(G1956), .B(G2474), .Z(new_n710));
  XOR2_X1   g285(.A(G1961), .B(G1966), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n709), .A2(new_n714), .A3(new_n712), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n717));
  AOI211_X1 g292(.A(new_n713), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(G1981), .B(G1986), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(G229));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n668), .B2(new_n730), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n735), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n734), .B1(new_n737), .B2(G1966), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G1966), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(G5), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G171), .B2(new_n735), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n739), .B1(G1961), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G34), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n730), .B1(new_n745), .B2(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(KEYINPUT98), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(KEYINPUT98), .B2(new_n747), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G160), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n730), .A2(G27), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT100), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n503), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2078), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n484), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(G129), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT26), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(G105), .B2(new_n656), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n730), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n730), .B2(G32), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n752), .B(new_n756), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n730), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n484), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n482), .A2(G128), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n470), .A2(G116), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n470), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n484), .A2(G139), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G33), .B(new_n786), .S(G29), .Z(new_n787));
  INV_X1    g362(.A(G1341), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n570), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G16), .B2(G19), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n787), .A2(G2072), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n769), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n767), .A2(new_n768), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n788), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n787), .A2(G2072), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  INV_X1    g372(.A(new_n741), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n743), .A2(new_n744), .A3(new_n792), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G2090), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT29), .Z(new_n804));
  AOI21_X1  g379(.A(new_n800), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n735), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1956), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n804), .B2(new_n801), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n735), .A2(G4), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n643), .B2(new_n735), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(KEYINPUT101), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n805), .A2(new_n811), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT33), .B(G1976), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n735), .A2(G23), .ZN(new_n819));
  INV_X1    g394(.A(G288), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n735), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(KEYINPUT92), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(KEYINPUT92), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n735), .A2(G6), .ZN(new_n825));
  INV_X1    g400(.A(G305), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n735), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT32), .B(G1981), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT91), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n822), .A2(new_n823), .A3(new_n818), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n735), .A2(G22), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT93), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G166), .B2(new_n735), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1971), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G1971), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n837), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT94), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n833), .A2(new_n834), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n845));
  MUX2_X1   g420(.A(G24), .B(G290), .S(G16), .Z(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT90), .B(G1986), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n484), .A2(G131), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n482), .A2(G119), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n470), .A2(G107), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  MUX2_X1   g428(.A(G25), .B(new_n853), .S(G29), .Z(new_n854));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G1991), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n848), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n844), .A2(new_n845), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n845), .B1(new_n844), .B2(new_n858), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n833), .A2(new_n840), .A3(new_n843), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT34), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n862), .B2(KEYINPUT34), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n860), .A2(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT36), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n859), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n817), .B1(new_n868), .B2(new_n873), .ZN(G311));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n868), .ZN(new_n875));
  INV_X1    g450(.A(new_n817), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(G150));
  NAND2_X1  g452(.A1(new_n536), .A2(G93), .ZN(new_n878));
  INV_X1    g453(.A(G55), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n562), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n531), .A2(G67), .A3(new_n533), .ZN(new_n881));
  NAND2_X1  g456(.A1(G80), .A2(G543), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n519), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G860), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n643), .A2(G559), .ZN(new_n888));
  XOR2_X1   g463(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n570), .A2(new_n884), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n566), .A2(new_n569), .B1(new_n880), .B2(new_n883), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n890), .B(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(KEYINPUT39), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n885), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n887), .B1(new_n895), .B2(new_n896), .ZN(G145));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n668), .B(new_n475), .ZN(new_n899));
  XNOR2_X1  g474(.A(G162), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n484), .A2(G142), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n482), .A2(G130), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n470), .A2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n658), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n853), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n776), .B(G164), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(new_n786), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n786), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(new_n764), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n764), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(new_n908), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n916), .A2(new_n917), .A3(new_n912), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n901), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n915), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n913), .A2(KEYINPUT103), .A3(new_n908), .A4(new_n914), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n900), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n918), .A2(KEYINPUT103), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n898), .B(new_n919), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(new_n893), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n651), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G299), .A2(new_n640), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n586), .B(new_n631), .C1(new_n638), .C2(new_n639), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n643), .A2(new_n649), .A3(new_n893), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n928), .A2(new_n932), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT41), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n926), .B(new_n933), .C1(new_n934), .C2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n928), .B2(new_n932), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n620), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n626), .B2(new_n623), .ZN(new_n944));
  INV_X1    g519(.A(new_n627), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n826), .ZN(new_n946));
  AOI21_X1  g521(.A(G305), .B1(new_n625), .B2(new_n627), .ZN(new_n947));
  AND3_X1   g522(.A1(G288), .A2(new_n528), .A3(new_n524), .ZN(new_n948));
  AOI21_X1  g523(.A(G288), .B1(new_n528), .B2(new_n524), .ZN(new_n949));
  OAI22_X1  g524(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G288), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n826), .B1(new_n944), .B2(new_n945), .ZN(new_n952));
  INV_X1    g527(.A(new_n524), .ZN(new_n953));
  INV_X1    g528(.A(new_n528), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n820), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n625), .A2(G305), .A3(new_n627), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n951), .A2(new_n952), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n939), .A2(new_n942), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n939), .B2(new_n942), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G868), .B2(new_n884), .ZN(G295));
  OAI21_X1  g538(.A(new_n962), .B1(G868), .B2(new_n884), .ZN(G331));
  INV_X1    g539(.A(new_n931), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n602), .A2(G171), .ZN(new_n966));
  NAND2_X1  g541(.A1(G301), .A2(new_n548), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(new_n893), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n893), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G301), .B1(new_n599), .B2(new_n601), .ZN(new_n971));
  NOR2_X1   g546(.A1(G171), .A2(G168), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n927), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n893), .A3(new_n967), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n936), .A3(new_n937), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n959), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n958), .A3(new_n975), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n970), .A2(new_n958), .A3(new_n975), .A4(KEYINPUT104), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n977), .A2(new_n980), .A3(new_n984), .A4(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n982), .A2(new_n989), .A3(KEYINPUT43), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n985), .B2(KEYINPUT105), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n976), .A2(new_n959), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n994), .A2(new_n898), .A3(new_n981), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n984), .A4(new_n980), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT107), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n988), .C1(new_n992), .C2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(G397));
  XNOR2_X1  g578(.A(new_n776), .B(new_n778), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n765), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n468), .B1(new_n472), .B2(G125), .ZN(new_n1007));
  OAI211_X1 g582(.A(G40), .B(new_n474), .C1(new_n1007), .C2(new_n470), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n469), .A2(KEYINPUT108), .A3(G40), .A4(new_n474), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n503), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT109), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n765), .A2(new_n1015), .A3(new_n1005), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n853), .A2(new_n856), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n853), .A2(new_n856), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G290), .A2(G1986), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT114), .B(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n503), .B2(new_n1013), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1012), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n503), .A2(new_n1031), .A3(new_n1013), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT111), .B(G2090), .Z(new_n1035));
  AND3_X1   g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1013), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1012), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G1971), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1030), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n1042));
  NAND4_X1  g617(.A1(G303), .A2(new_n1042), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n524), .A2(new_n528), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT113), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n524), .A2(G8), .A3(new_n528), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT112), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1043), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1028), .B(new_n1041), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1045), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1044), .A2(KEYINPUT113), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1052), .A2(new_n1053), .B1(new_n1054), .B2(KEYINPUT112), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1034), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n503), .A2(KEYINPUT110), .A3(new_n1031), .A4(new_n1013), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n841), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1056), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1043), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1055), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1029), .B1(new_n1064), .B2(new_n1014), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n820), .A2(G1976), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G305), .A2(G1981), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G305), .A2(G1981), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1077), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n1070), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(new_n1071), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1073), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1051), .A2(new_n1069), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1055), .A2(new_n1068), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1028), .B1(new_n1087), .B2(new_n1041), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1010), .B(new_n1011), .C1(new_n1014), .C2(new_n1031), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n797), .B1(new_n1092), .B2(new_n1060), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT119), .A4(new_n443), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT53), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT119), .B1(new_n1039), .B2(new_n443), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1091), .B(new_n1093), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1065), .B2(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1065), .B2(G2078), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(KEYINPUT53), .A3(new_n1094), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1091), .B1(new_n1103), .B2(new_n1093), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1090), .B(G171), .C1(new_n1100), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT120), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1099), .A3(new_n1097), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1090), .B1(new_n1109), .B2(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1089), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1061), .A2(KEYINPUT116), .A3(new_n1033), .A4(new_n751), .ZN(new_n1113));
  INV_X1    g688(.A(G1966), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1065), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1092), .A2(new_n1060), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT116), .B1(new_n1117), .B2(new_n751), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n548), .A2(new_n1030), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1112), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n548), .B(new_n1030), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1118), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1030), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT51), .B1(new_n548), .B2(new_n1030), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1121), .A2(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1027), .B1(new_n1111), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT51), .A3(new_n1122), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(G171), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1105), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(new_n1139), .A3(KEYINPUT123), .A4(new_n1089), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT124), .B1(new_n1128), .B2(KEYINPUT62), .ZN(new_n1141));
  AND4_X1   g716(.A1(KEYINPUT124), .A2(new_n1132), .A3(KEYINPUT62), .A4(new_n1133), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1130), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1087), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n1085), .A3(new_n1067), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1081), .A2(new_n1082), .A3(new_n820), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1070), .B1(new_n1147), .B2(new_n1077), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1087), .A2(new_n1041), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT115), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1069), .A2(new_n1085), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n1051), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1125), .A2(new_n602), .A3(new_n1030), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1150), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(new_n1153), .C1(new_n1145), .C2(new_n1067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1149), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1008), .A2(new_n1098), .A3(G2078), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1063), .A2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT122), .Z(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n1093), .A3(new_n1099), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1164), .A2(G171), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT54), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1167));
  INV_X1    g742(.A(G1956), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n586), .B(KEYINPUT57), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(new_n442), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1039), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1012), .A2(G1384), .A3(G164), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT58), .B(G1341), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1065), .A2(G1996), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1180), .B2(new_n570), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1180), .A2(new_n570), .ZN(new_n1182));
  AND2_X1   g757(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n814), .B1(new_n1092), .B2(new_n1060), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1178), .A2(new_n778), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT60), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n642), .A3(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1190), .A2(new_n642), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1176), .A2(new_n1184), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1170), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1187), .A2(new_n642), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1174), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1164), .A2(G171), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1198), .B(KEYINPUT54), .C1(new_n1109), .C2(G171), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1197), .A2(new_n1128), .A3(new_n1089), .A4(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1159), .B1(new_n1166), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1026), .B1(new_n1144), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1017), .A2(new_n1019), .A3(new_n1018), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(G2067), .B2(new_n776), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1016), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1015), .A2(new_n1005), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT46), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n1004), .A2(new_n765), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n1210), .B2(new_n1016), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1211), .B(new_n1212), .Z(new_n1213));
  NAND3_X1  g788(.A1(new_n1204), .A2(KEYINPUT125), .A3(new_n1016), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1024), .A2(new_n1015), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT48), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1022), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1207), .A2(new_n1213), .A3(new_n1214), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1218), .B(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1202), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g796(.A1(G227), .A2(new_n461), .ZN(new_n1223));
  OAI21_X1  g797(.A(new_n1223), .B1(new_n726), .B2(new_n727), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n691), .B2(new_n692), .ZN(new_n1225));
  NAND3_X1  g799(.A1(new_n1225), .A2(new_n924), .A3(new_n986), .ZN(G225));
  INV_X1    g800(.A(G225), .ZN(G308));
endmodule


