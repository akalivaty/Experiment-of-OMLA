

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808;

  XOR2_X1 U374 ( .A(KEYINPUT9), .B(G122), .Z(n560) );
  XNOR2_X1 U375 ( .A(G143), .B(G122), .ZN(n547) );
  XNOR2_X1 U376 ( .A(KEYINPUT16), .B(G122), .ZN(n570) );
  INV_X1 U377 ( .A(G146), .ZN(n591) );
  AND2_X2 U378 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X2 U379 ( .A(n618), .B(n379), .ZN(n635) );
  NOR2_X2 U380 ( .A1(n609), .A2(n608), .ZN(n357) );
  XOR2_X2 U381 ( .A(n533), .B(n532), .Z(n375) );
  AND2_X2 U382 ( .A1(n480), .A2(n372), .ZN(n478) );
  XNOR2_X2 U383 ( .A(n602), .B(n601), .ZN(n646) );
  XNOR2_X2 U384 ( .A(n352), .B(KEYINPUT109), .ZN(n630) );
  NAND2_X2 U385 ( .A1(n473), .A2(n698), .ZN(n352) );
  XNOR2_X1 U386 ( .A(G119), .B(G110), .ZN(n526) );
  XNOR2_X1 U387 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n549) );
  XNOR2_X1 U388 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n573) );
  INV_X1 U389 ( .A(G237), .ZN(n582) );
  NAND2_X1 U390 ( .A1(n623), .A2(n622), .ZN(n734) );
  BUF_X1 U391 ( .A(n466), .Z(n463) );
  BUF_X1 U392 ( .A(G953), .Z(n443) );
  BUF_X1 U393 ( .A(G116), .Z(n449) );
  BUF_X1 U394 ( .A(G128), .Z(n447) );
  BUF_X1 U395 ( .A(G107), .Z(n450) );
  AND2_X1 U396 ( .A1(n480), .A2(n483), .ZN(n353) );
  AND2_X2 U397 ( .A1(n440), .A2(n438), .ZN(n437) );
  NOR2_X2 U398 ( .A1(n688), .A2(n784), .ZN(n689) );
  XNOR2_X1 U399 ( .A(n362), .B(KEYINPUT85), .ZN(n637) );
  XNOR2_X2 U400 ( .A(n566), .B(n576), .ZN(n587) );
  XNOR2_X2 U401 ( .A(n577), .B(G134), .ZN(n566) );
  NOR2_X2 U402 ( .A1(n719), .A2(n736), .ZN(n606) );
  INV_X1 U403 ( .A(n721), .ZN(n698) );
  NOR2_X2 U404 ( .A1(G953), .A2(G237), .ZN(n545) );
  AND2_X1 U405 ( .A1(n423), .A2(n422), .ZN(n421) );
  OR2_X1 U406 ( .A1(n467), .A2(G902), .ZN(n520) );
  NAND2_X1 U407 ( .A1(G237), .A2(G234), .ZN(n355) );
  XNOR2_X2 U408 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U409 ( .A1(n507), .A2(n506), .ZN(n365) );
  AND2_X1 U410 ( .A1(n504), .A2(n386), .ZN(n503) );
  AND2_X1 U411 ( .A1(n476), .A2(n491), .ZN(n490) );
  NAND2_X1 U412 ( .A1(n408), .A2(n458), .ZN(n407) );
  NAND2_X1 U413 ( .A1(n436), .A2(KEYINPUT36), .ZN(n435) );
  NAND2_X1 U414 ( .A1(n460), .A2(n376), .ZN(n404) );
  XNOR2_X1 U415 ( .A(n462), .B(n461), .ZN(n460) );
  XNOR2_X1 U416 ( .A(n357), .B(KEYINPUT76), .ZN(n453) );
  XNOR2_X1 U417 ( .A(n605), .B(KEYINPUT103), .ZN(n736) );
  NAND2_X2 U418 ( .A1(n401), .A2(n398), .ZN(n607) );
  INV_X1 U419 ( .A(n371), .ZN(n354) );
  AND2_X1 U420 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U421 ( .A(n704), .B(KEYINPUT59), .ZN(n705) );
  XNOR2_X1 U422 ( .A(n528), .B(n511), .ZN(n529) );
  XNOR2_X1 U423 ( .A(n469), .B(G146), .ZN(n468) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n536) );
  XNOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .ZN(n581) );
  XNOR2_X1 U426 ( .A(G131), .B(G140), .ZN(n586) );
  XNOR2_X1 U427 ( .A(G131), .B(KEYINPUT5), .ZN(n516) );
  XNOR2_X1 U428 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n356) );
  AND2_X2 U429 ( .A1(n417), .A2(n679), .ZN(n680) );
  NAND2_X1 U430 ( .A1(n681), .A2(n680), .ZN(n476) );
  NAND2_X1 U431 ( .A1(n637), .A2(n731), .ZN(n762) );
  NAND2_X1 U432 ( .A1(n359), .A2(n358), .ZN(n609) );
  INV_X1 U433 ( .A(n607), .ZN(n358) );
  INV_X1 U434 ( .A(n638), .ZN(n359) );
  NOR2_X1 U435 ( .A1(n388), .A2(n581), .ZN(n491) );
  NAND2_X1 U436 ( .A1(n360), .A2(n405), .ZN(n369) );
  NAND2_X1 U437 ( .A1(n406), .A2(n724), .ZN(n360) );
  NAND2_X1 U438 ( .A1(n370), .A2(n367), .ZN(n366) );
  AND2_X2 U439 ( .A1(n466), .A2(n749), .ZN(n659) );
  XNOR2_X2 U440 ( .A(n361), .B(n486), .ZN(n775) );
  NAND2_X1 U441 ( .A1(n487), .A2(n490), .ZN(n361) );
  NAND2_X1 U442 ( .A1(n363), .A2(n634), .ZN(n362) );
  XNOR2_X1 U443 ( .A(n364), .B(n492), .ZN(n363) );
  NAND2_X1 U444 ( .A1(n494), .A2(n493), .ZN(n364) );
  NAND2_X1 U445 ( .A1(n365), .A2(n386), .ZN(n502) );
  NOR2_X1 U446 ( .A1(n365), .A2(n706), .ZN(n497) );
  AND2_X1 U447 ( .A1(n659), .A2(n354), .ZN(n639) );
  XNOR2_X2 U448 ( .A(n366), .B(n412), .ZN(n411) );
  INV_X1 U449 ( .A(n707), .ZN(n368) );
  NAND2_X1 U450 ( .A1(n700), .A2(KEYINPUT44), .ZN(n370) );
  XNOR2_X2 U451 ( .A(n404), .B(KEYINPUT35), .ZN(n700) );
  XNOR2_X1 U452 ( .A(n520), .B(n519), .ZN(n371) );
  XNOR2_X1 U453 ( .A(n520), .B(n519), .ZN(n668) );
  OR2_X1 U454 ( .A1(n778), .A2(n399), .ZN(n398) );
  XNOR2_X2 U455 ( .A(n607), .B(n597), .ZN(n466) );
  NAND2_X1 U456 ( .A1(n805), .A2(n713), .ZN(n672) );
  XNOR2_X1 U457 ( .A(n456), .B(n556), .ZN(n704) );
  NAND2_X1 U458 ( .A1(n672), .A2(KEYINPUT44), .ZN(n477) );
  INV_X1 U459 ( .A(n736), .ZN(n405) );
  NAND2_X1 U460 ( .A1(n774), .A2(G902), .ZN(n402) );
  AND2_X1 U461 ( .A1(n675), .A2(n416), .ZN(n415) );
  NAND2_X1 U462 ( .A1(n672), .A2(n413), .ZN(n416) );
  XNOR2_X1 U463 ( .A(n446), .B(n445), .ZN(n561) );
  INV_X1 U464 ( .A(KEYINPUT8), .ZN(n445) );
  NAND2_X1 U465 ( .A1(n785), .A2(G234), .ZN(n446) );
  NOR2_X1 U466 ( .A1(n417), .A2(KEYINPUT2), .ZN(n388) );
  NAND2_X1 U467 ( .A1(n488), .A2(n763), .ZN(n487) );
  INV_X1 U468 ( .A(KEYINPUT75), .ZN(n489) );
  XNOR2_X1 U469 ( .A(n660), .B(KEYINPUT33), .ZN(n739) );
  XNOR2_X1 U470 ( .A(n568), .B(n567), .ZN(n623) );
  INV_X1 U471 ( .A(KEYINPUT1), .ZN(n597) );
  INV_X1 U472 ( .A(G137), .ZN(n469) );
  XNOR2_X1 U473 ( .A(n471), .B(n516), .ZN(n470) );
  XNOR2_X1 U474 ( .A(n449), .B(n450), .ZN(n559) );
  OR2_X1 U475 ( .A1(n705), .A2(n702), .ZN(n505) );
  NAND2_X1 U476 ( .A1(n784), .A2(n508), .ZN(n501) );
  INV_X1 U477 ( .A(n431), .ZN(n430) );
  NAND2_X1 U478 ( .A1(n426), .A2(n382), .ZN(n423) );
  NAND2_X1 U479 ( .A1(n374), .A2(n433), .ZN(n425) );
  AND2_X1 U480 ( .A1(n431), .A2(n381), .ZN(n420) );
  INV_X1 U481 ( .A(KEYINPUT123), .ZN(n429) );
  INV_X1 U482 ( .A(KEYINPUT48), .ZN(n492) );
  INV_X1 U483 ( .A(n744), .ZN(n510) );
  NOR2_X1 U484 ( .A1(KEYINPUT87), .A2(n414), .ZN(n413) );
  INV_X1 U485 ( .A(KEYINPUT44), .ZN(n414) );
  INV_X1 U486 ( .A(KEYINPUT88), .ZN(n412) );
  XNOR2_X1 U487 ( .A(G137), .B(KEYINPUT68), .ZN(n593) );
  XNOR2_X1 U488 ( .A(G113), .B(G104), .ZN(n553) );
  INV_X1 U489 ( .A(KEYINPUT10), .ZN(n522) );
  XOR2_X1 U490 ( .A(KEYINPUT79), .B(KEYINPUT23), .Z(n524) );
  XNOR2_X1 U491 ( .A(n447), .B(G140), .ZN(n523) );
  XNOR2_X1 U492 ( .A(n454), .B(n527), .ZN(n528) );
  XNOR2_X1 U493 ( .A(n526), .B(n455), .ZN(n454) );
  INV_X1 U494 ( .A(KEYINPUT24), .ZN(n455) );
  NAND2_X1 U495 ( .A1(n682), .A2(n583), .ZN(n483) );
  NAND2_X1 U496 ( .A1(n581), .A2(n482), .ZN(n481) );
  INV_X1 U497 ( .A(n583), .ZN(n482) );
  XNOR2_X1 U498 ( .A(n558), .B(n457), .ZN(n622) );
  XNOR2_X1 U499 ( .A(n557), .B(n702), .ZN(n457) );
  NAND2_X1 U500 ( .A1(G469), .A2(n400), .ZN(n399) );
  INV_X1 U501 ( .A(KEYINPUT105), .ZN(n651) );
  XNOR2_X1 U502 ( .A(n668), .B(n377), .ZN(n658) );
  INV_X1 U503 ( .A(KEYINPUT65), .ZN(n486) );
  OR2_X1 U504 ( .A1(n434), .A2(G469), .ZN(n432) );
  NAND2_X1 U505 ( .A1(n661), .A2(n739), .ZN(n462) );
  INV_X1 U506 ( .A(KEYINPUT34), .ZN(n461) );
  XNOR2_X1 U507 ( .A(n470), .B(n468), .ZN(n517) );
  XNOR2_X1 U508 ( .A(n564), .B(n444), .ZN(n782) );
  XOR2_X1 U509 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n563) );
  AND2_X1 U510 ( .A1(n463), .A2(n439), .ZN(n438) );
  NAND2_X1 U511 ( .A1(n391), .A2(KEYINPUT36), .ZN(n439) );
  XNOR2_X1 U512 ( .A(n667), .B(n452), .ZN(n805) );
  INV_X1 U513 ( .A(KEYINPUT32), .ZN(n452) );
  NAND2_X1 U514 ( .A1(n465), .A2(n464), .ZN(n657) );
  INV_X1 U515 ( .A(n743), .ZN(n464) );
  INV_X1 U516 ( .A(n504), .ZN(n498) );
  NAND2_X1 U517 ( .A1(n420), .A2(n424), .ZN(n419) );
  NAND2_X1 U518 ( .A1(n428), .A2(n427), .ZN(n424) );
  AND2_X1 U519 ( .A1(n483), .A2(n479), .ZN(n372) );
  XOR2_X1 U520 ( .A(n778), .B(n777), .Z(n373) );
  AND2_X1 U521 ( .A1(n432), .A2(n485), .ZN(n374) );
  XOR2_X1 U522 ( .A(n663), .B(n662), .Z(n376) );
  XOR2_X1 U523 ( .A(n521), .B(KEYINPUT6), .Z(n377) );
  NOR2_X1 U524 ( .A1(n463), .A2(n629), .ZN(n378) );
  INV_X1 U525 ( .A(G902), .ZN(n400) );
  XNOR2_X1 U526 ( .A(KEYINPUT39), .B(KEYINPUT72), .ZN(n379) );
  XOR2_X1 U527 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n380) );
  INV_X1 U528 ( .A(KEYINPUT36), .ZN(n495) );
  INV_X1 U529 ( .A(n433), .ZN(n427) );
  NAND2_X1 U530 ( .A1(n434), .A2(G469), .ZN(n433) );
  AND2_X1 U531 ( .A1(n374), .A2(n429), .ZN(n381) );
  AND2_X1 U532 ( .A1(n425), .A2(KEYINPUT123), .ZN(n382) );
  INV_X1 U533 ( .A(G469), .ZN(n774) );
  XOR2_X1 U534 ( .A(n467), .B(KEYINPUT62), .Z(n383) );
  XNOR2_X1 U535 ( .A(KEYINPUT86), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U536 ( .A(n394), .B(KEYINPUT124), .Z(n385) );
  INV_X1 U537 ( .A(KEYINPUT87), .ZN(n458) );
  INV_X1 U538 ( .A(n373), .ZN(n434) );
  INV_X1 U539 ( .A(n706), .ZN(n508) );
  AND2_X1 U540 ( .A1(n485), .A2(n706), .ZN(n386) );
  XNOR2_X1 U541 ( .A(n534), .B(n375), .ZN(n387) );
  XNOR2_X1 U542 ( .A(n534), .B(n375), .ZN(n543) );
  BUF_X2 U543 ( .A(n775), .Z(n703) );
  NAND2_X1 U544 ( .A1(n703), .A2(n374), .ZN(n426) );
  NAND2_X1 U545 ( .A1(n703), .A2(n705), .ZN(n507) );
  INV_X1 U546 ( .A(n609), .ZN(n389) );
  OR2_X1 U547 ( .A1(n417), .A2(KEYINPUT2), .ZN(n390) );
  BUF_X1 U548 ( .A(n602), .Z(n391) );
  NAND2_X1 U549 ( .A1(n437), .A2(n435), .ZN(n392) );
  NAND2_X1 U550 ( .A1(n437), .A2(n435), .ZN(n729) );
  XNOR2_X2 U551 ( .A(n795), .B(n596), .ZN(n778) );
  XNOR2_X1 U552 ( .A(n396), .B(KEYINPUT94), .ZN(n406) );
  XNOR2_X1 U553 ( .A(n650), .B(KEYINPUT93), .ZN(n397) );
  NAND2_X1 U554 ( .A1(n397), .A2(n371), .ZN(n396) );
  BUF_X1 U555 ( .A(n635), .Z(n393) );
  BUF_X1 U556 ( .A(n693), .Z(n394) );
  BUF_X1 U557 ( .A(n630), .Z(n395) );
  INV_X1 U558 ( .A(n406), .ZN(n697) );
  NAND2_X1 U559 ( .A1(n778), .A2(n774), .ZN(n403) );
  NAND2_X2 U560 ( .A1(n409), .A2(n407), .ZN(n677) );
  INV_X1 U561 ( .A(n411), .ZN(n408) );
  AND2_X2 U562 ( .A1(n410), .A2(n415), .ZN(n409) );
  NAND2_X1 U563 ( .A1(n411), .A2(n459), .ZN(n410) );
  NAND2_X1 U564 ( .A1(n417), .A2(n785), .ZN(n789) );
  XNOR2_X2 U565 ( .A(n677), .B(n676), .ZN(n417) );
  XNOR2_X1 U566 ( .A(n762), .B(n489), .ZN(n488) );
  NOR2_X2 U567 ( .A1(n806), .A2(n808), .ZN(n628) );
  XNOR2_X2 U568 ( .A(n418), .B(n593), .ZN(n796) );
  XNOR2_X1 U569 ( .A(n418), .B(n546), .ZN(n556) );
  XNOR2_X2 U570 ( .A(n575), .B(n522), .ZN(n418) );
  INV_X1 U571 ( .A(n703), .ZN(n428) );
  NAND2_X1 U572 ( .A1(n421), .A2(n419), .ZN(G54) );
  NAND2_X1 U573 ( .A1(n430), .A2(KEYINPUT123), .ZN(n422) );
  NAND2_X1 U574 ( .A1(n703), .A2(n373), .ZN(n431) );
  NAND2_X1 U575 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U576 ( .A(n630), .B(KEYINPUT112), .ZN(n442) );
  INV_X1 U577 ( .A(n442), .ZN(n436) );
  AND2_X1 U578 ( .A1(n585), .A2(n495), .ZN(n441) );
  INV_X2 U579 ( .A(G125), .ZN(n509) );
  XNOR2_X2 U580 ( .A(n513), .B(n512), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n566), .B(n565), .ZN(n444) );
  INV_X1 U582 ( .A(n784), .ZN(n485) );
  NAND2_X1 U583 ( .A1(n478), .A2(n484), .ZN(n602) );
  XNOR2_X2 U584 ( .A(n571), .B(n448), .ZN(n790) );
  XNOR2_X2 U585 ( .A(n590), .B(n570), .ZN(n448) );
  XNOR2_X2 U586 ( .A(n515), .B(n514), .ZN(n571) );
  NAND2_X1 U587 ( .A1(n635), .A2(n698), .ZN(n620) );
  INV_X1 U588 ( .A(n658), .ZN(n656) );
  NAND2_X1 U589 ( .A1(n598), .A2(n658), .ZN(n475) );
  XNOR2_X2 U590 ( .A(n612), .B(KEYINPUT38), .ZN(n732) );
  XNOR2_X2 U591 ( .A(n451), .B(n624), .ZN(n767) );
  NOR2_X2 U592 ( .A1(n735), .A2(n734), .ZN(n451) );
  XNOR2_X2 U593 ( .A(n796), .B(n525), .ZN(n530) );
  XNOR2_X2 U594 ( .A(n790), .B(n580), .ZN(n684) );
  AND2_X2 U595 ( .A1(n453), .A2(n611), .ZN(n617) );
  XNOR2_X2 U596 ( .A(n530), .B(n529), .ZN(n693) );
  XNOR2_X1 U597 ( .A(n628), .B(n384), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n555), .B(n554), .ZN(n456) );
  AND2_X1 U599 ( .A1(n477), .A2(KEYINPUT87), .ZN(n459) );
  NAND2_X1 U600 ( .A1(n463), .A2(n743), .ZN(n664) );
  INV_X1 U601 ( .A(n463), .ZN(n465) );
  NOR2_X1 U602 ( .A1(n669), .A2(n463), .ZN(n670) );
  NOR2_X1 U603 ( .A1(n749), .A2(n463), .ZN(n750) );
  XNOR2_X1 U604 ( .A(n587), .B(n518), .ZN(n467) );
  NAND2_X1 U605 ( .A1(n545), .A2(G210), .ZN(n471) );
  XNOR2_X1 U606 ( .A(n475), .B(n474), .ZN(n473) );
  INV_X1 U607 ( .A(KEYINPUT108), .ZN(n474) );
  AND2_X1 U608 ( .A1(n476), .A2(n390), .ZN(n765) );
  OR2_X2 U609 ( .A1(n684), .A2(n481), .ZN(n480) );
  NAND2_X1 U610 ( .A1(n484), .A2(n353), .ZN(n612) );
  INV_X1 U611 ( .A(n629), .ZN(n479) );
  NAND2_X1 U612 ( .A1(n684), .A2(n583), .ZN(n484) );
  XNOR2_X2 U613 ( .A(n587), .B(n586), .ZN(n795) );
  INV_X2 U614 ( .A(n775), .ZN(n779) );
  XNOR2_X1 U615 ( .A(n616), .B(KEYINPUT69), .ZN(n494) );
  NAND2_X1 U616 ( .A1(n499), .A2(n496), .ZN(G60) );
  NAND2_X1 U617 ( .A1(n498), .A2(n497), .ZN(n496) );
  NOR2_X1 U618 ( .A1(n503), .A2(n500), .ZN(n499) );
  NAND2_X1 U619 ( .A1(n502), .A2(n501), .ZN(n500) );
  NOR2_X1 U620 ( .A1(n703), .A2(n505), .ZN(n504) );
  NAND2_X1 U621 ( .A1(n705), .A2(n702), .ZN(n506) );
  XNOR2_X2 U622 ( .A(n509), .B(G146), .ZN(n575) );
  INV_X1 U623 ( .A(n387), .ZN(n743) );
  NAND2_X1 U624 ( .A1(n387), .A2(n510), .ZN(n638) );
  NOR2_X2 U625 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X2 U626 ( .A1(n693), .A2(G902), .ZN(n534) );
  AND2_X1 U627 ( .A1(n561), .A2(G221), .ZN(n511) );
  INV_X1 U628 ( .A(n701), .ZN(n634) );
  BUF_X1 U629 ( .A(n739), .Z(n766) );
  XNOR2_X2 U630 ( .A(G143), .B(G128), .ZN(n577) );
  XNOR2_X2 U631 ( .A(G101), .B(G116), .ZN(n513) );
  XNOR2_X2 U632 ( .A(G113), .B(KEYINPUT71), .ZN(n512) );
  XNOR2_X1 U633 ( .A(KEYINPUT3), .B(G119), .ZN(n514) );
  XNOR2_X1 U634 ( .A(n517), .B(n571), .ZN(n518) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(G472), .ZN(n519) );
  INV_X1 U636 ( .A(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U637 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U638 ( .A(KEYINPUT83), .B(KEYINPUT92), .Z(n527) );
  INV_X4 U639 ( .A(G953), .ZN(n785) );
  XOR2_X1 U640 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n533) );
  NAND2_X1 U641 ( .A1(G234), .A2(n581), .ZN(n531) );
  XNOR2_X1 U642 ( .A(KEYINPUT20), .B(n531), .ZN(n540) );
  NAND2_X1 U643 ( .A1(n540), .A2(G217), .ZN(n532) );
  NAND2_X1 U644 ( .A1(n536), .A2(G952), .ZN(n535) );
  XOR2_X1 U645 ( .A(KEYINPUT89), .B(n535), .Z(n761) );
  NOR2_X1 U646 ( .A1(n443), .A2(n761), .ZN(n643) );
  NAND2_X1 U647 ( .A1(G902), .A2(n536), .ZN(n641) );
  NOR2_X1 U648 ( .A1(G900), .A2(n641), .ZN(n537) );
  NAND2_X1 U649 ( .A1(n443), .A2(n537), .ZN(n538) );
  XNOR2_X1 U650 ( .A(KEYINPUT107), .B(n538), .ZN(n539) );
  NOR2_X1 U651 ( .A1(n643), .A2(n539), .ZN(n608) );
  NAND2_X1 U652 ( .A1(n540), .A2(G221), .ZN(n541) );
  XNOR2_X1 U653 ( .A(n541), .B(KEYINPUT21), .ZN(n744) );
  OR2_X1 U654 ( .A1(n608), .A2(n744), .ZN(n542) );
  XNOR2_X1 U655 ( .A(n544), .B(KEYINPUT70), .ZN(n598) );
  NAND2_X1 U656 ( .A1(G214), .A2(n545), .ZN(n546) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n548) );
  XNOR2_X1 U658 ( .A(n548), .B(n547), .ZN(n552) );
  XOR2_X1 U659 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n550) );
  XNOR2_X1 U660 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U661 ( .A(n552), .B(n551), .ZN(n555) );
  XOR2_X1 U662 ( .A(n553), .B(n586), .Z(n554) );
  NOR2_X1 U663 ( .A1(G902), .A2(n704), .ZN(n558) );
  XNOR2_X1 U664 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n557) );
  INV_X1 U665 ( .A(G475), .ZN(n702) );
  XNOR2_X1 U666 ( .A(n560), .B(n559), .ZN(n565) );
  NAND2_X1 U667 ( .A1(G217), .A2(n561), .ZN(n562) );
  XNOR2_X1 U668 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U669 ( .A1(n782), .A2(n400), .ZN(n568) );
  XOR2_X1 U670 ( .A(KEYINPUT102), .B(G478), .Z(n567) );
  INV_X1 U671 ( .A(n623), .ZN(n604) );
  OR2_X1 U672 ( .A1(n622), .A2(n604), .ZN(n721) );
  XNOR2_X2 U673 ( .A(G110), .B(G107), .ZN(n569) );
  XNOR2_X2 U674 ( .A(n569), .B(G104), .ZN(n590) );
  NAND2_X1 U675 ( .A1(n785), .A2(G224), .ZN(n572) );
  XNOR2_X1 U676 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U677 ( .A(n575), .B(n574), .ZN(n579) );
  XNOR2_X1 U678 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U679 ( .A(n579), .B(n578), .ZN(n580) );
  INV_X1 U680 ( .A(n581), .ZN(n682) );
  NAND2_X1 U681 ( .A1(n400), .A2(n582), .ZN(n584) );
  NAND2_X1 U682 ( .A1(n584), .A2(G210), .ZN(n583) );
  AND2_X1 U683 ( .A1(n584), .A2(G214), .ZN(n629) );
  INV_X1 U684 ( .A(n391), .ZN(n585) );
  NAND2_X1 U685 ( .A1(n785), .A2(G227), .ZN(n588) );
  XNOR2_X1 U686 ( .A(n588), .B(KEYINPUT80), .ZN(n589) );
  XNOR2_X1 U687 ( .A(n590), .B(n589), .ZN(n595) );
  XNOR2_X1 U688 ( .A(n591), .B(G101), .ZN(n592) );
  XNOR2_X1 U689 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U690 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U691 ( .A1(n598), .A2(n354), .ZN(n599) );
  XNOR2_X1 U692 ( .A(n599), .B(KEYINPUT28), .ZN(n600) );
  NOR2_X1 U693 ( .A1(n600), .A2(n607), .ZN(n625) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n601) );
  INV_X1 U695 ( .A(n646), .ZN(n603) );
  NAND2_X1 U696 ( .A1(n625), .A2(n603), .ZN(n719) );
  NAND2_X1 U697 ( .A1(n622), .A2(n604), .ZN(n725) );
  NAND2_X1 U698 ( .A1(n721), .A2(n725), .ZN(n605) );
  XNOR2_X1 U699 ( .A(n606), .B(KEYINPUT47), .ZN(n614) );
  NOR2_X1 U700 ( .A1(n371), .A2(n629), .ZN(n610) );
  XNOR2_X1 U701 ( .A(KEYINPUT30), .B(n610), .ZN(n611) );
  OR2_X1 U702 ( .A1(n622), .A2(n623), .ZN(n663) );
  NOR2_X1 U703 ( .A1(n663), .A2(n612), .ZN(n613) );
  NAND2_X1 U704 ( .A1(n617), .A2(n613), .ZN(n718) );
  AND2_X1 U705 ( .A1(n614), .A2(n718), .ZN(n615) );
  NAND2_X1 U706 ( .A1(n729), .A2(n615), .ZN(n616) );
  NAND2_X1 U707 ( .A1(n617), .A2(n732), .ZN(n618) );
  INV_X1 U708 ( .A(KEYINPUT40), .ZN(n619) );
  XNOR2_X1 U709 ( .A(n620), .B(n619), .ZN(n806) );
  NAND2_X1 U710 ( .A1(n732), .A2(n479), .ZN(n621) );
  XNOR2_X1 U711 ( .A(n621), .B(KEYINPUT110), .ZN(n735) );
  XNOR2_X1 U712 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n767), .A2(n625), .ZN(n627) );
  INV_X1 U714 ( .A(KEYINPUT42), .ZN(n626) );
  XNOR2_X1 U715 ( .A(n627), .B(n626), .ZN(n808) );
  NAND2_X1 U716 ( .A1(n395), .A2(n378), .ZN(n631) );
  XOR2_X1 U717 ( .A(KEYINPUT43), .B(n631), .Z(n633) );
  INV_X1 U718 ( .A(n612), .ZN(n632) );
  NOR2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n701) );
  INV_X1 U720 ( .A(n725), .ZN(n709) );
  NAND2_X1 U721 ( .A1(n393), .A2(n709), .ZN(n731) );
  NAND2_X1 U722 ( .A1(n731), .A2(KEYINPUT2), .ZN(n678) );
  NAND2_X1 U723 ( .A1(n678), .A2(KEYINPUT82), .ZN(n636) );
  AND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n681) );
  INV_X1 U725 ( .A(n638), .ZN(n749) );
  XNOR2_X1 U726 ( .A(n639), .B(KEYINPUT95), .ZN(n753) );
  NOR2_X1 U727 ( .A1(G898), .A2(n785), .ZN(n640) );
  XOR2_X1 U728 ( .A(KEYINPUT90), .B(n640), .Z(n791) );
  NOR2_X1 U729 ( .A1(n791), .A2(n641), .ZN(n642) );
  OR2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U731 ( .A(n644), .B(KEYINPUT91), .ZN(n645) );
  NOR2_X2 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X2 U733 ( .A(n647), .B(n380), .ZN(n661) );
  INV_X1 U734 ( .A(n661), .ZN(n648) );
  NOR2_X1 U735 ( .A1(n753), .A2(n648), .ZN(n649) );
  XNOR2_X1 U736 ( .A(n649), .B(KEYINPUT31), .ZN(n724) );
  NAND2_X1 U737 ( .A1(n661), .A2(n389), .ZN(n650) );
  NOR2_X1 U738 ( .A1(n744), .A2(n734), .ZN(n652) );
  XNOR2_X1 U739 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U740 ( .A1(n653), .A2(n661), .ZN(n655) );
  INV_X1 U741 ( .A(KEYINPUT22), .ZN(n654) );
  XNOR2_X2 U742 ( .A(n655), .B(n654), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(n656), .ZN(n666) );
  NOR2_X1 U744 ( .A1(n666), .A2(n657), .ZN(n707) );
  NAND2_X1 U745 ( .A1(n659), .A2(n658), .ZN(n660) );
  INV_X1 U746 ( .A(KEYINPUT81), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n664), .B(KEYINPUT106), .ZN(n665) );
  NOR2_X1 U748 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n743), .A2(n371), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n713) );
  INV_X1 U751 ( .A(n672), .ZN(n674) );
  NOR2_X1 U752 ( .A1(n700), .A2(KEYINPUT44), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U754 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n676) );
  OR2_X1 U755 ( .A1(n678), .A2(KEYINPUT82), .ZN(n679) );
  INV_X1 U756 ( .A(KEYINPUT2), .ZN(n763) );
  NAND2_X1 U757 ( .A1(n779), .A2(G210), .ZN(n686) );
  XOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n683) );
  XNOR2_X1 U759 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n686), .B(n685), .ZN(n688) );
  INV_X1 U761 ( .A(G952), .ZN(n687) );
  AND2_X1 U762 ( .A1(n687), .A2(n443), .ZN(n784) );
  XNOR2_X1 U763 ( .A(n689), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U764 ( .A1(n779), .A2(G472), .ZN(n690) );
  XNOR2_X1 U765 ( .A(n690), .B(n383), .ZN(n691) );
  NAND2_X1 U766 ( .A1(n691), .A2(n485), .ZN(n692) );
  XNOR2_X1 U767 ( .A(n692), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U768 ( .A1(n779), .A2(G217), .ZN(n694) );
  XNOR2_X1 U769 ( .A(n694), .B(n385), .ZN(n695) );
  NAND2_X1 U770 ( .A1(n695), .A2(n485), .ZN(n696) );
  XNOR2_X1 U771 ( .A(n696), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n697), .A2(n698), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n699), .B(G104), .ZN(G6) );
  XOR2_X1 U774 ( .A(n700), .B(G122), .Z(G24) );
  XOR2_X1 U775 ( .A(G140), .B(n701), .Z(G42) );
  XNOR2_X1 U776 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n706) );
  XNOR2_X1 U777 ( .A(G101), .B(n707), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n708), .B(KEYINPUT113), .ZN(G3) );
  XNOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n697), .A2(n709), .ZN(n710) );
  XOR2_X1 U781 ( .A(n711), .B(n710), .Z(n712) );
  XNOR2_X1 U782 ( .A(n450), .B(n712), .ZN(G9) );
  XNOR2_X1 U783 ( .A(G110), .B(KEYINPUT114), .ZN(n714) );
  XNOR2_X1 U784 ( .A(n714), .B(n713), .ZN(G12) );
  NOR2_X1 U785 ( .A1(n719), .A2(n725), .ZN(n716) );
  XNOR2_X1 U786 ( .A(n447), .B(KEYINPUT29), .ZN(n715) );
  XNOR2_X1 U787 ( .A(n716), .B(n715), .ZN(G30) );
  XOR2_X1 U788 ( .A(G143), .B(KEYINPUT115), .Z(n717) );
  XNOR2_X1 U789 ( .A(n718), .B(n717), .ZN(G45) );
  NOR2_X1 U790 ( .A1(n719), .A2(n721), .ZN(n720) );
  XOR2_X1 U791 ( .A(G146), .B(n720), .Z(G48) );
  NOR2_X1 U792 ( .A1(n721), .A2(n724), .ZN(n722) );
  XOR2_X1 U793 ( .A(KEYINPUT116), .B(n722), .Z(n723) );
  XNOR2_X1 U794 ( .A(G113), .B(n723), .ZN(G15) );
  NOR2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U796 ( .A(n449), .B(KEYINPUT117), .ZN(n726) );
  XNOR2_X1 U797 ( .A(n727), .B(n726), .ZN(G18) );
  XOR2_X1 U798 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n728) );
  XNOR2_X1 U799 ( .A(n392), .B(n728), .ZN(n730) );
  XNOR2_X1 U800 ( .A(G125), .B(n730), .ZN(G27) );
  XNOR2_X1 U801 ( .A(G134), .B(n731), .ZN(G36) );
  NOR2_X1 U802 ( .A1(n732), .A2(n479), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U804 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n741) );
  INV_X1 U806 ( .A(n766), .ZN(n740) );
  NOR2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U808 ( .A(n742), .B(KEYINPUT121), .ZN(n758) );
  XOR2_X1 U809 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n746) );
  NAND2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U811 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U812 ( .A(n747), .B(KEYINPUT119), .ZN(n748) );
  NOR2_X1 U813 ( .A1(n748), .A2(n354), .ZN(n752) );
  XOR2_X1 U814 ( .A(KEYINPUT50), .B(n750), .Z(n751) );
  NAND2_X1 U815 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U816 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U817 ( .A(KEYINPUT51), .B(n755), .Z(n756) );
  NAND2_X1 U818 ( .A1(n756), .A2(n767), .ZN(n757) );
  NAND2_X1 U819 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U820 ( .A(KEYINPUT52), .B(n759), .Z(n760) );
  NOR2_X1 U821 ( .A1(n761), .A2(n760), .ZN(n771) );
  BUF_X1 U822 ( .A(n762), .Z(n797) );
  NAND2_X1 U823 ( .A1(n797), .A2(n763), .ZN(n764) );
  NAND2_X1 U824 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U825 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U826 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U827 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U828 ( .A1(n785), .A2(n772), .ZN(n773) );
  XOR2_X1 U829 ( .A(KEYINPUT53), .B(n773), .Z(G75) );
  XNOR2_X1 U830 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n776) );
  XNOR2_X1 U831 ( .A(n776), .B(KEYINPUT57), .ZN(n777) );
  BUF_X1 U832 ( .A(n779), .Z(n780) );
  NAND2_X1 U833 ( .A1(n780), .A2(G478), .ZN(n781) );
  XOR2_X1 U834 ( .A(n782), .B(n781), .Z(n783) );
  NOR2_X1 U835 ( .A1(n784), .A2(n783), .ZN(G63) );
  NAND2_X1 U836 ( .A1(n443), .A2(G224), .ZN(n786) );
  XNOR2_X1 U837 ( .A(KEYINPUT61), .B(n786), .ZN(n787) );
  NAND2_X1 U838 ( .A1(n787), .A2(G898), .ZN(n788) );
  NAND2_X1 U839 ( .A1(n789), .A2(n788), .ZN(n794) );
  XNOR2_X1 U840 ( .A(n790), .B(KEYINPUT126), .ZN(n792) );
  NAND2_X1 U841 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U842 ( .A(n794), .B(n793), .Z(G69) );
  XNOR2_X1 U843 ( .A(n796), .B(n795), .ZN(n800) );
  XNOR2_X1 U844 ( .A(n797), .B(n800), .ZN(n798) );
  NOR2_X1 U845 ( .A1(n798), .A2(n443), .ZN(n799) );
  XNOR2_X1 U846 ( .A(n799), .B(KEYINPUT127), .ZN(n804) );
  XOR2_X1 U847 ( .A(G227), .B(n800), .Z(n801) );
  NAND2_X1 U848 ( .A1(n801), .A2(G900), .ZN(n802) );
  NAND2_X1 U849 ( .A1(n802), .A2(n443), .ZN(n803) );
  NAND2_X1 U850 ( .A1(n804), .A2(n803), .ZN(G72) );
  XNOR2_X1 U851 ( .A(n805), .B(G119), .ZN(G21) );
  BUF_X1 U852 ( .A(n806), .Z(n807) );
  XOR2_X1 U853 ( .A(G131), .B(n807), .Z(G33) );
  XOR2_X1 U854 ( .A(n808), .B(G137), .Z(G39) );
endmodule

