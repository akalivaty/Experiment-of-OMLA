//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n202), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G226gat), .A2(G233gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n216), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n230));
  AND4_X1   g029(.A1(new_n224), .A2(new_n227), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(G183gat), .B(G190gat), .C1(KEYINPUT66), .C2(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n222), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n233), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n245), .A3(new_n241), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n222), .A4(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n223), .B2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n229), .A3(KEYINPUT27), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n227), .A4(new_n230), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT27), .B(G183gat), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT26), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n220), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n219), .B2(KEYINPUT71), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n218), .A2(new_n262), .A3(new_n259), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n233), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n238), .B(new_n247), .C1(new_n258), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n215), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n222), .A2(new_n244), .A3(new_n246), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n269), .A2(new_n243), .B1(new_n237), .B2(KEYINPUT25), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n264), .A2(new_n233), .ZN(new_n271));
  INV_X1    g070(.A(new_n255), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n227), .A2(new_n230), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT67), .B(G183gat), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(KEYINPUT27), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n275), .B2(new_n252), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n257), .A2(new_n256), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n214), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n213), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n266), .A2(new_n215), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT29), .B1(new_n270), .B2(new_n278), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n281), .B(new_n212), .C1(new_n282), .C2(new_n215), .ZN(new_n283));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT78), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n280), .A2(new_n283), .A3(new_n290), .A4(new_n287), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT37), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n293), .A3(new_n283), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n286), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n280), .B2(new_n283), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT38), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G57gat), .B(G85gat), .Z(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G1gat), .B(G29gat), .Z(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT84), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n300), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(KEYINPUT72), .B2(new_n314), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n312), .A2(G120gat), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n306), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n305), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n310), .A2(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(KEYINPUT2), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G155gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n330));
  OAI21_X1  g129(.A(G162gat), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n324), .B1(new_n331), .B2(KEYINPUT2), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(G141gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n322), .A2(KEYINPUT82), .A3(new_n326), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  INV_X1    g139(.A(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n327), .A2(G155gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n323), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n326), .B1(new_n346), .B2(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n320), .A2(new_n321), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n318), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n314), .B2(new_n313), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(new_n309), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n340), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n347), .A2(new_n351), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(KEYINPUT4), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(KEYINPUT81), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n348), .B(new_n361), .C1(new_n350), .C2(new_n309), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n326), .C1(new_n346), .C2(new_n336), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(new_n360), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n354), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n360), .A2(new_n347), .A3(new_n362), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n339), .A3(new_n352), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n356), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n369), .A3(KEYINPUT5), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n353), .B1(new_n347), .B2(new_n351), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n353), .B1(new_n339), .B2(new_n352), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n304), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n370), .A2(new_n376), .A3(new_n304), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT6), .B(new_n304), .C1(new_n370), .C2(new_n376), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n292), .B(new_n297), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n283), .A2(KEYINPUT92), .ZN(new_n384));
  INV_X1    g183(.A(new_n268), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n281), .A4(new_n212), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n387), .A3(new_n280), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT37), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT38), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n294), .A2(new_n390), .A3(new_n286), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT93), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT93), .B1(new_n389), .B2(new_n391), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n364), .A2(new_n267), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n213), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n210), .B2(new_n211), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n347), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n212), .B1(new_n364), .B2(new_n267), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n399), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n396), .B(new_n398), .C1(KEYINPUT86), .C2(new_n400), .ZN(new_n405));
  AOI21_X1  g204(.A(G22gat), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(G22gat), .A3(new_n405), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n401), .B1(new_n403), .B2(new_n402), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n398), .B2(new_n396), .ZN(new_n412));
  INV_X1    g211(.A(new_n405), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n407), .B(new_n410), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(new_n406), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n408), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n419), .A2(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT88), .B1(new_n409), .B2(new_n418), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n383), .A2(new_n394), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n289), .A2(new_n427), .A3(new_n291), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n287), .B1(new_n280), .B2(new_n283), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n280), .A2(new_n283), .A3(new_n287), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(KEYINPUT30), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n428), .A2(KEYINPUT90), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT90), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n365), .A2(new_n371), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n435), .B(new_n356), .C1(new_n436), .C2(new_n373), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n355), .B1(new_n372), .B2(new_n374), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n367), .A2(new_n339), .A3(new_n355), .A4(new_n352), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n304), .B(new_n437), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n377), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n356), .B1(new_n436), .B2(new_n373), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT39), .A3(new_n439), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(KEYINPUT40), .A3(new_n304), .A4(new_n437), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT91), .B1(new_n434), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n451));
  NOR4_X1   g250(.A1(new_n432), .A2(new_n433), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n426), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT94), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n431), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n428), .A2(new_n431), .A3(KEYINPUT90), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n451), .B1(new_n459), .B2(new_n448), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n434), .A2(KEYINPUT91), .A3(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n426), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n266), .A2(new_n322), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT64), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n270), .A2(new_n278), .A3(new_n351), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT32), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT74), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n476), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n469), .B(KEYINPUT32), .C1(new_n471), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n465), .A2(new_n468), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT75), .B(KEYINPUT34), .C1(new_n481), .C2(new_n467), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT75), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n467), .B1(new_n465), .B2(new_n468), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n480), .A2(new_n488), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n480), .B(new_n488), .Z(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n419), .A2(new_n420), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n423), .A2(new_n421), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n425), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n379), .A2(new_n378), .ZN(new_n501));
  OR3_X1    g300(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n377), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n377), .B1(new_n501), .B2(KEYINPUT85), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n455), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n494), .B1(new_n495), .B2(new_n497), .C1(new_n500), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n495), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n493), .B1(new_n508), .B2(new_n496), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT89), .C1(new_n504), .C2(new_n500), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n454), .A2(new_n464), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n500), .A2(new_n495), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n380), .A2(new_n381), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n459), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT11), .ZN(new_n522));
  INV_X1    g321(.A(G169gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(G197gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G1gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  MUX2_X1   g328(.A(G1gat), .B(new_n528), .S(new_n529), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G8gat), .ZN(new_n531));
  NOR3_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(KEYINPUT95), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(KEYINPUT95), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G43gat), .B(G50gat), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(KEYINPUT96), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n534), .A2(new_n535), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n539), .A2(KEYINPUT97), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n540), .ZN(new_n550));
  INV_X1    g349(.A(new_n532), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n551), .A2(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n531), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n547), .A2(new_n557), .A3(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n559), .B2(new_n531), .ZN(new_n560));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n555), .B(new_n531), .Z(new_n563));
  XOR2_X1   g362(.A(new_n561), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT18), .B1(new_n560), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n526), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  INV_X1    g368(.A(new_n526), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n562), .A3(new_n565), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n520), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT103), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT101), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n576), .B2(KEYINPUT7), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT101), .A3(G85gat), .A4(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n583), .A3(KEYINPUT7), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n575), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n575), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n558), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n557), .B1(new_n547), .B2(new_n553), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n559), .A2(KEYINPUT102), .A3(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n593), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n555), .A2(new_n601), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n600), .B2(new_n603), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n574), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n600), .A2(new_n603), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n604), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT103), .A3(new_n606), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n609), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n615), .A2(KEYINPUT103), .A3(new_n606), .A4(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620));
  INV_X1    g419(.A(G64gat), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(G57gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n621), .A2(G57gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(new_n626), .B2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT9), .B1(new_n622), .B2(new_n624), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n628), .A3(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n531), .B1(new_n637), .B2(new_n636), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n646), .B2(new_n651), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n620), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  INV_X1    g455(.A(new_n620), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n619), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n619), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n593), .A2(new_n636), .ZN(new_n664));
  INV_X1    g463(.A(new_n636), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n592), .A3(new_n591), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n664), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n665), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT105), .B1(new_n674), .B2(new_n668), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n676), .B(new_n669), .C1(new_n672), .C2(new_n673), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n670), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n668), .ZN(new_n683));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n670), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n661), .A2(new_n663), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n573), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n502), .A2(new_n503), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT106), .B(G1gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1324gat));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n434), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT16), .B(G8gat), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT107), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(G8gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT107), .B(new_n700), .C1(new_n695), .C2(new_n696), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(G1325gat));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n689), .A2(new_n703), .A3(new_n495), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n573), .A2(new_n509), .A3(new_n688), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n703), .ZN(G1326gat));
  INV_X1    g505(.A(new_n500), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NAND2_X1  g509(.A1(new_n655), .A2(new_n658), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n687), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n619), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n520), .A2(new_n572), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n690), .A2(G29gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n617), .A2(new_n618), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n511), .B2(new_n519), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n572), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n568), .A2(new_n571), .A3(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n712), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n505), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n453), .A2(KEYINPUT94), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n463), .B1(new_n462), .B2(new_n426), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n514), .A2(new_n515), .B1(new_n512), .B2(new_n517), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n619), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n720), .B(new_n725), .C1(new_n731), .C2(KEYINPUT44), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n732), .B2(new_n690), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n733), .A3(new_n734), .ZN(G1328gat));
  NOR3_X1   g534(.A1(new_n714), .A2(G36gat), .A3(new_n459), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n732), .B2(new_n459), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n714), .A2(new_n508), .ZN(new_n740));
  INV_X1    g539(.A(new_n509), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n740), .A2(G43gat), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n732), .A2(new_n746), .A3(new_n500), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n732), .B2(new_n500), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n714), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n520), .A2(KEYINPUT110), .A3(new_n572), .A4(new_n713), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n500), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT48), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n732), .A2(new_n500), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n753), .A2(new_n754), .B1(new_n757), .B2(G50gat), .ZN(new_n758));
  OAI22_X1  g557(.A1(new_n749), .A2(new_n756), .B1(new_n758), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n729), .A2(new_n730), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n661), .A2(new_n663), .A3(new_n686), .A4(new_n724), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n690), .B(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n434), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n768), .B2(new_n767), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n763), .A2(G71gat), .A3(new_n741), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n762), .A2(new_n508), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(G71gat), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n763), .A2(new_n707), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g576(.A1(new_n724), .A2(new_n711), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n731), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n505), .B1(new_n454), .B2(new_n464), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n718), .B(new_n780), .C1(new_n782), .C2(new_n519), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n691), .A2(new_n587), .A3(new_n686), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n780), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n687), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n720), .C1(new_n731), .C2(KEYINPUT44), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n690), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(G1336gat));
  OAI21_X1  g593(.A(G92gat), .B1(new_n792), .B2(new_n459), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT115), .B(G92gat), .C1(new_n792), .C2(new_n459), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n784), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n459), .A2(G92gat), .A3(new_n687), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n799), .A3(KEYINPUT51), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n797), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n786), .B2(new_n802), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n795), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  NOR3_X1   g608(.A1(new_n508), .A2(G99gat), .A3(new_n687), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n792), .B2(new_n509), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  NOR3_X1   g612(.A1(new_n500), .A2(G106gat), .A3(new_n687), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n801), .A2(new_n803), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n817), .A3(new_n803), .A4(new_n814), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n792), .B2(new_n500), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n786), .B2(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1339gat));
  NOR3_X1   g623(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT54), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n674), .B2(new_n668), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n672), .A2(new_n669), .A3(new_n673), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n684), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  INV_X1    g631(.A(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n834), .A3(new_n685), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT118), .A4(new_n685), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(new_n722), .A3(new_n723), .A4(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n525), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n560), .A2(new_n561), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n563), .A2(new_n564), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n571), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n686), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n718), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n617), .A2(new_n618), .A3(new_n844), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n711), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n661), .A2(new_n663), .A3(new_n687), .A4(new_n724), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n707), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n434), .A2(new_n690), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n495), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n572), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n312), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n850), .A2(new_n851), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n764), .A2(new_n459), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n512), .ZN(new_n860));
  INV_X1    g659(.A(new_n724), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n856), .B1(new_n862), .B2(new_n312), .ZN(G1340gat));
  NOR3_X1   g662(.A1(new_n854), .A2(new_n318), .A3(new_n687), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n686), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n318), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n867), .A3(new_n659), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n854), .B2(new_n711), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  INV_X1    g669(.A(new_n512), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(G134gat), .A3(new_n619), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n854), .B2(new_n619), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n741), .A2(new_n500), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n855), .A2(G141gat), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n857), .A2(new_n858), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n509), .A2(new_n853), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n500), .B1(new_n850), .B2(new_n851), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n572), .A2(new_n685), .A3(new_n831), .A4(new_n834), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n887), .A2(new_n845), .B1(new_n617), .B2(new_n618), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n711), .B1(new_n849), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n886), .B(new_n500), .C1(new_n851), .C2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n572), .B(new_n883), .C1(new_n885), .C2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n335), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n881), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n883), .B1(new_n885), .B2(new_n890), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n892), .B1(new_n897), .B2(new_n724), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n879), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n895), .A2(new_n896), .B1(new_n899), .B2(new_n880), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n500), .A2(KEYINPUT57), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n661), .A2(new_n855), .A3(new_n663), .A4(new_n687), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n848), .A2(new_n835), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n711), .B1(new_n904), .B2(new_n888), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n857), .A2(new_n707), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n686), .A3(new_n883), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G148gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT59), .ZN(new_n911));
  INV_X1    g710(.A(G148gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(KEYINPUT59), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n897), .B2(new_n687), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT120), .B(new_n913), .C1(new_n897), .C2(new_n687), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n859), .A2(new_n877), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n912), .A3(new_n686), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  OAI22_X1  g720(.A1(new_n897), .A2(new_n711), .B1(new_n328), .B2(new_n330), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n919), .A2(new_n342), .A3(new_n343), .A4(new_n659), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n897), .B2(new_n619), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n341), .A3(new_n718), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  OR2_X1    g726(.A1(new_n764), .A2(new_n459), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n508), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n852), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n523), .A3(new_n855), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n857), .A2(new_n690), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT121), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n871), .A2(new_n459), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n861), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n936), .B2(new_n523), .ZN(G1348gat));
  INV_X1    g736(.A(G176gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n938), .A3(new_n686), .ZN(new_n939));
  OAI21_X1  g738(.A(G176gat), .B1(new_n930), .B2(new_n687), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  NOR2_X1   g740(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n942));
  AND2_X1   g741(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n659), .A2(new_n256), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n934), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n274), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n930), .B2(new_n711), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n942), .B(new_n943), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  AND4_X1   g749(.A1(KEYINPUT122), .A2(new_n947), .A3(KEYINPUT60), .A4(new_n949), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1350gat));
  NOR2_X1   g751(.A1(new_n619), .A2(new_n273), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n934), .B(new_n953), .C1(new_n945), .C2(new_n946), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n852), .A2(new_n718), .A3(new_n929), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G190gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(new_n957), .A3(G190gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n956), .B1(new_n961), .B2(new_n963), .ZN(G1351gat));
  NOR2_X1   g763(.A1(new_n928), .A2(new_n741), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n908), .A2(KEYINPUT125), .A3(new_n572), .A4(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n903), .A2(new_n905), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n901), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n969), .B(new_n965), .C1(new_n884), .C2(new_n886), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n855), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n971), .A3(G197gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n877), .A2(new_n434), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n724), .A2(G197gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n933), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n972), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1352gat));
  NOR2_X1   g780(.A1(new_n687), .A2(G204gat), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n974), .B(new_n982), .C1(new_n945), .C2(new_n946), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n908), .A2(new_n686), .A3(new_n965), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n983), .A2(KEYINPUT62), .B1(new_n984), .B2(G204gat), .ZN(new_n985));
  INV_X1    g784(.A(new_n983), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT127), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n983), .A2(new_n989), .A3(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n985), .B1(new_n988), .B2(new_n990), .ZN(G1353gat));
  OAI21_X1  g790(.A(G211gat), .B1(new_n970), .B2(new_n711), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT63), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n933), .A2(new_n974), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n659), .A2(new_n205), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n970), .B2(new_n619), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n718), .A2(new_n206), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n995), .B2(new_n999), .ZN(G1355gat));
endmodule


