//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(KEYINPUT64), .A2(G113), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT64), .B1(G113), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n467), .A3(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n470), .A2(new_n476), .A3(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT66), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G124), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n483), .A2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n462), .A2(new_n465), .A3(new_n467), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n474), .A2(new_n467), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n488), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(G543), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(new_n516), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n508), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n511), .A2(new_n532), .B1(new_n533), .B2(new_n516), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n525), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n506), .A2(new_n510), .A3(G81), .ZN(new_n540));
  OAI211_X1 g115(.A(G43), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n540), .A2(KEYINPUT68), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT68), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(KEYINPUT69), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n525), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n510), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  OR2_X1    g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n504), .A2(new_n505), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n567), .B2(G91), .ZN(new_n568));
  AND4_X1   g143(.A1(new_n564), .A2(new_n506), .A3(new_n510), .A4(G91), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n558), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n572));
  XNOR2_X1  g147(.A(G168), .B(new_n572), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n525), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  INV_X1    g152(.A(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n565), .B2(new_n566), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n567), .B2(G87), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n567), .A2(new_n582), .A3(G87), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n525), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n567), .B2(G86), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n579), .A2(new_n592), .A3(G48), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT74), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n525), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n508), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(new_n600), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n567), .A2(G85), .B1(new_n579), .B2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n511), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n516), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n525), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n614), .A2(new_n615), .B1(new_n618), .B2(G651), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n606), .B1(G868), .B2(new_n620), .ZN(G284));
  OAI21_X1  g196(.A(new_n606), .B1(G868), .B2(new_n620), .ZN(G321));
  NOR2_X1   g197(.A1(G299), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G286), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  AOI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n611), .A2(new_n619), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g209(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n638), .A2(new_n639), .B1(KEYINPUT77), .B2(G2100), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  NOR2_X1   g216(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n488), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n481), .B2(G135), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n649), .ZN(G156));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT80), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(KEYINPUT80), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n655), .A2(G2427), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G2427), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n653), .A2(KEYINPUT80), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(new_n654), .ZN(new_n660));
  OAI21_X1  g235(.A(G2430), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT79), .B(G2438), .Z(new_n662));
  OAI21_X1  g237(.A(G2427), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  INV_X1    g238(.A(G2430), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n658), .A3(new_n654), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT14), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n662), .B1(new_n661), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n652), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n661), .A2(new_n666), .ZN(new_n674));
  INV_X1    g249(.A(new_n662), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n652), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n676), .A2(KEYINPUT14), .A3(new_n667), .A4(new_n677), .ZN(new_n678));
  AND3_X1   g253(.A1(new_n670), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n673), .B1(new_n670), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1341), .B(G1348), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT81), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n651), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n670), .A2(new_n678), .ZN(new_n686));
  INV_X1    g261(.A(new_n673), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n670), .A2(new_n673), .A3(new_n678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n683), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n685), .B(new_n691), .C1(new_n679), .C2(new_n680), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n684), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G401));
  XNOR2_X1  g271(.A(G2084), .B(G2090), .ZN(new_n697));
  XNOR2_X1  g272(.A(G2067), .B(G2678), .ZN(new_n698));
  XNOR2_X1  g273(.A(G2072), .B(G2078), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(KEYINPUT17), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n698), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT83), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(new_n697), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT18), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n698), .A2(new_n697), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n703), .B(new_n706), .C1(new_n701), .C2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G2096), .B(G2100), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(G227));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1971), .B(G1976), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1956), .B(G2474), .Z(new_n716));
  XOR2_X1   g291(.A(G1961), .B(G1966), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n716), .A2(new_n717), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(new_n718), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n721), .B1(new_n715), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n715), .A2(new_n722), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT20), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(G1991), .B(G1996), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n728), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n724), .B2(new_n726), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n731), .B1(new_n729), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n712), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n729), .A2(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(new_n730), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(new_n711), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(G229));
  NAND3_X1  g316(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT25), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n495), .A2(G127), .ZN(new_n744));
  INV_X1    g319(.A(G115), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n464), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n743), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n481), .A2(G139), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n751), .B2(G33), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n751), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n751), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n648), .A2(G29), .ZN(new_n760));
  AND2_X1   g335(.A1(KEYINPUT30), .A2(G28), .ZN(new_n761));
  NOR2_X1   g336(.A1(KEYINPUT30), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n751), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G11), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(new_n751), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  INV_X1    g343(.A(G160), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n751), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n772), .B1(new_n771), .B2(new_n770), .C1(new_n753), .C2(new_n754), .ZN(new_n773));
  INV_X1    g348(.A(G16), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n756), .A2(new_n759), .A3(new_n773), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n774), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n774), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1961), .ZN(new_n783));
  NOR2_X1   g358(.A1(G168), .A2(new_n774), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n774), .B2(G21), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n786), .B2(G1966), .ZN(new_n787));
  INV_X1    g362(.A(G1966), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(new_n788), .B1(G1961), .B2(new_n782), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT26), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n792), .A2(new_n793), .B1(new_n477), .B2(G105), .ZN(new_n794));
  INV_X1    g369(.A(G129), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n488), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n481), .B2(G141), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n751), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n751), .B2(G32), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n787), .B(new_n789), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n751), .A2(G26), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT28), .Z(new_n803));
  NAND3_X1  g378(.A1(new_n489), .A2(KEYINPUT94), .A3(G128), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n805));
  INV_X1    g380(.A(G128), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n488), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(G116), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(G2105), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n481), .B2(G140), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n803), .B1(new_n813), .B2(G29), .ZN(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n774), .A2(G4), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n620), .B2(new_n774), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1348), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n801), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n780), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n548), .A2(new_n774), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n774), .B2(G19), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT93), .B(G1341), .Z(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n799), .A2(new_n800), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT97), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n751), .A2(G35), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G162), .B2(new_n751), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT29), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G2090), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n821), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n774), .A2(G23), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n586), .B2(new_n774), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G1976), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(KEYINPUT33), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G1976), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n774), .A2(G22), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G166), .B2(new_n774), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT91), .Z(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(G1971), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(G1971), .ZN(new_n850));
  MUX2_X1   g425(.A(G6), .B(G305), .S(G16), .Z(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT32), .B(G1981), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n843), .A2(new_n845), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT34), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G1991), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n751), .A2(G25), .ZN(new_n859));
  OR2_X1    g434(.A1(G95), .A2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n861));
  INV_X1    g436(.A(G119), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n488), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G131), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n468), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT85), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT86), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n859), .B1(new_n870), .B2(G29), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT87), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n855), .A2(new_n856), .B1(new_n858), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n858), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n774), .A2(G24), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT88), .Z(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(G290), .B2(G16), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT89), .B(G1986), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n843), .A2(new_n845), .A3(new_n854), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT34), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n873), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT36), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT92), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n873), .A2(new_n887), .A3(new_n880), .A4(new_n882), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n835), .B1(new_n886), .B2(new_n888), .ZN(G311));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n834), .ZN(G150));
  XNOR2_X1  g466(.A(KEYINPUT98), .B(G93), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n567), .A2(new_n892), .B1(new_n579), .B2(G55), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n508), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n893), .B(KEYINPUT99), .C1(new_n508), .C2(new_n894), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G860), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n620), .A2(G559), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT101), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n546), .A2(new_n547), .A3(new_n895), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n544), .A3(new_n898), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(KEYINPUT100), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n905), .B(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n913), .A2(KEYINPUT39), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n900), .B1(new_n913), .B2(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n902), .B1(new_n914), .B2(new_n915), .ZN(G145));
  XNOR2_X1  g491(.A(new_n769), .B(new_n648), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(G162), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n797), .A2(new_n812), .A3(new_n808), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n797), .B1(new_n808), .B2(new_n812), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n750), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n502), .B(KEYINPUT102), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n797), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n813), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n749), .A3(new_n919), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  OR2_X1    g505(.A1(G106), .A2(G2105), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n932));
  INV_X1    g507(.A(G130), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n488), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G142), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n468), .A2(new_n935), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n934), .A2(new_n936), .A3(new_n637), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n637), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n867), .A2(new_n937), .A3(new_n868), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n938), .A2(new_n937), .B1(new_n867), .B2(new_n868), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n930), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n869), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(KEYINPUT103), .A3(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n924), .B1(new_n922), .B2(new_n927), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n929), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n922), .A2(new_n927), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n923), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n950), .A2(new_n928), .B1(new_n945), .B2(new_n942), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n918), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n929), .B2(new_n947), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n928), .A3(new_n939), .A4(new_n944), .ZN(new_n955));
  INV_X1    g530(.A(new_n918), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g534(.A(KEYINPUT106), .B1(new_n899), .B2(G868), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(G303), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n586), .B(G305), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n961), .B(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n912), .A2(new_n630), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n910), .A2(new_n631), .A3(new_n911), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n968));
  NAND2_X1  g543(.A1(G299), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G91), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT71), .B1(new_n511), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n567), .A2(new_n564), .A3(G91), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(KEYINPUT104), .A3(new_n563), .A4(new_n558), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n620), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n629), .A2(new_n968), .A3(G299), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT41), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n979), .B(new_n980), .C1(new_n975), .C2(new_n976), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n975), .A2(new_n980), .A3(new_n976), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n975), .B2(new_n976), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n984), .B2(new_n979), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n966), .A3(new_n965), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n964), .A2(new_n978), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G868), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n964), .B1(new_n978), .B2(new_n986), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  MUX2_X1   g565(.A(new_n960), .B(KEYINPUT106), .S(new_n990), .Z(G295));
  MUX2_X1   g566(.A(new_n960), .B(KEYINPUT106), .S(new_n990), .Z(G331));
  NOR2_X1   g567(.A1(G171), .A2(G168), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G286), .B2(G301), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n906), .A2(KEYINPUT100), .A3(new_n907), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT100), .B1(new_n906), .B2(new_n907), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n910), .A2(new_n911), .A3(new_n995), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n985), .ZN(new_n1002));
  INV_X1    g577(.A(new_n963), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1000), .A3(new_n977), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1005), .A2(new_n953), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n999), .A2(new_n1000), .A3(new_n977), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n984), .B1(new_n999), .B2(new_n1000), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT107), .B(new_n963), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n963), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND4_X1   g587(.A1(KEYINPUT43), .A2(new_n1006), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1005), .A2(new_n953), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT44), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1006), .A2(new_n1019), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT43), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1018), .B1(KEYINPUT44), .B2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n497), .B2(new_n501), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1027));
  NOR2_X1   g602(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n497), .B2(new_n501), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G40), .A3(G160), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1027), .A2(new_n1030), .A3(G2084), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n473), .A2(new_n475), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G2105), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n465), .A2(new_n467), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(G137), .A3(new_n466), .A4(new_n462), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1035), .A3(G40), .A4(new_n478), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G1384), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n502), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1026), .A2(new_n1037), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1031), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G166), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT55), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(G1971), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1036), .B1(new_n502), .B2(new_n1028), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1044), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1043), .B(KEYINPUT63), .C1(new_n1046), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n591), .A2(new_n596), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1057), .A2(KEYINPUT117), .A3(KEYINPUT49), .A4(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1026), .A2(new_n1036), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1044), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT49), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT116), .B(KEYINPUT49), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1064), .B(new_n1066), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1054), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1048), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1046), .B(G8), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n842), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n577), .A2(new_n580), .ZN(new_n1077));
  INV_X1    g652(.A(new_n585), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(G1976), .C1(new_n1078), .C2(new_n583), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1075), .A2(new_n1076), .A3(new_n1066), .A4(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(G8), .C1(new_n1026), .C2(new_n1036), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n586), .B2(G1976), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(KEYINPUT52), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1071), .A2(new_n1074), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1056), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1046), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1036), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1053), .A2(new_n1090), .A3(new_n1029), .ZN(new_n1091));
  AOI21_X1  g666(.A(G2090), .B1(new_n1091), .B2(KEYINPUT118), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1051), .A2(new_n1093), .A3(new_n1053), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1073), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT119), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1095), .B2(KEYINPUT119), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1089), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1087), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1043), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1052), .A3(new_n1094), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1050), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(G8), .A3(new_n1096), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1087), .B1(new_n1110), .B2(new_n1089), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1101), .B1(new_n1111), .B2(new_n1043), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1088), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1071), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1074), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1071), .A2(new_n842), .A3(new_n586), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1059), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1066), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1961), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1091), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G2078), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1039), .A2(KEYINPUT53), .A3(new_n1121), .A4(new_n1040), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1047), .B2(G2078), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G168), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G8), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1042), .A2(KEYINPUT51), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1040), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1038), .B1(new_n497), .B2(new_n501), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1090), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n788), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1051), .A2(new_n771), .A3(new_n1053), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1130), .B(G8), .C1(new_n1136), .C2(new_n1127), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1128), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT124), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1140), .B(new_n1128), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1129), .B(new_n1137), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1126), .B1(new_n1142), .B2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1142), .B2(KEYINPUT62), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1144), .A3(KEYINPUT62), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT57), .ZN(new_n1148));
  XNOR2_X1  g723(.A(G299), .B(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1091), .A2(new_n778), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT56), .B(G2072), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1039), .A2(new_n1040), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1026), .A2(new_n1036), .A3(G2067), .ZN(new_n1154));
  INV_X1    g729(.A(G1348), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1091), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n629), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1150), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1156), .A2(KEYINPUT60), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT123), .B(new_n629), .C1(new_n1156), .C2(KEYINPUT60), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1155), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1154), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1165), .B2(new_n620), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n629), .A4(new_n1164), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT122), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1160), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1158), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(new_n1153), .A3(KEYINPUT61), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1149), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1176), .B2(new_n1158), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(G1341), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1047), .A2(G1996), .B1(new_n1065), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT59), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n548), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1180), .B2(new_n548), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1172), .A2(new_n1177), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1159), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1137), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1125), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(G171), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT54), .B1(new_n1190), .B2(new_n1126), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(G171), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT54), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1123), .A2(G301), .A3(new_n1125), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1129), .A2(new_n1188), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1146), .A2(new_n1147), .B1(new_n1185), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1111), .B(KEYINPUT125), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1113), .B(new_n1118), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1040), .A2(KEYINPUT108), .A3(new_n1036), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT108), .B1(new_n1040), .B2(new_n1036), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(G290), .A2(G1986), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT109), .ZN(new_n1205));
  AND2_X1   g780(.A1(G290), .A2(G1986), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1203), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT113), .ZN(new_n1208));
  INV_X1    g783(.A(G1996), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1203), .A2(new_n1209), .A3(new_n797), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT110), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1202), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1200), .A2(KEYINPUT110), .A3(new_n1201), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n797), .A2(new_n1209), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1215), .A2(KEYINPUT111), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1215), .A2(KEYINPUT111), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n813), .A2(G2067), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n808), .A2(new_n815), .A3(new_n812), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1212), .A2(new_n1213), .A3(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT112), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1208), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT112), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1222), .B(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1215), .B(KEYINPUT111), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1226), .A2(new_n1227), .A3(KEYINPUT113), .A4(new_n1210), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n869), .B(new_n858), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AND4_X1   g806(.A1(new_n1207), .A2(new_n1224), .A3(new_n1228), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1199), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1229), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n870), .A2(new_n858), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1224), .A2(new_n1228), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1234), .B1(new_n1236), .B2(new_n1220), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT48), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1224), .A2(new_n1228), .A3(new_n1231), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1203), .A2(new_n1209), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(KEYINPUT46), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1229), .B1(new_n925), .B2(new_n1221), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1244), .B(KEYINPUT47), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g821(.A1(new_n1237), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1233), .A2(new_n1247), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g823(.A1(G227), .A2(new_n459), .ZN(new_n1250));
  AOI21_X1  g824(.A(new_n1250), .B1(new_n736), .B2(new_n740), .ZN(new_n1251));
  NAND3_X1  g825(.A1(new_n695), .A2(new_n1251), .A3(new_n958), .ZN(new_n1252));
  INV_X1    g826(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g827(.A(KEYINPUT127), .B1(new_n1022), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1255));
  AOI211_X1 g829(.A(new_n1255), .B(new_n1252), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1256));
  NOR2_X1   g830(.A1(new_n1254), .A2(new_n1256), .ZN(G308));
  NAND2_X1  g831(.A1(new_n1022), .A2(new_n1253), .ZN(G225));
endmodule


