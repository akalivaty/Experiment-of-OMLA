//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT23), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n204), .A2(KEYINPUT65), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT65), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G183gat), .B(G190gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n210), .B(new_n212), .C1(new_n213), .C2(new_n209), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT25), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n202), .A2(new_n203), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT26), .B1(new_n202), .B2(new_n203), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n205), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  AOI21_X1  g022(.A(G190gat), .B1(new_n223), .B2(KEYINPUT27), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n225), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT28), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n212), .A3(new_n205), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n234), .B1(new_n237), .B2(KEYINPUT24), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n204), .A2(new_n212), .A3(new_n240), .A4(new_n205), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n233), .A2(new_n238), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n215), .A2(new_n231), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n248), .A2(new_n249), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n253), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n249), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT34), .ZN(new_n261));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n254), .A2(new_n258), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n215), .A2(new_n231), .A3(new_n263), .A4(new_n242), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT34), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n260), .B2(new_n264), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT32), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n271), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n270), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n262), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n238), .B(new_n212), .C1(new_n207), .C2(new_n206), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n239), .B(new_n210), .C1(new_n213), .C2(new_n209), .ZN(new_n286));
  AND4_X1   g085(.A1(new_n240), .A2(new_n204), .A3(new_n212), .A4(new_n205), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(KEYINPUT25), .A2(new_n285), .B1(new_n288), .B2(new_n233), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n263), .B1(new_n289), .B2(new_n231), .ZN(new_n290));
  INV_X1    g089(.A(new_n264), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n284), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n278), .B1(new_n292), .B2(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n279), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n277), .B1(new_n271), .B2(new_n272), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n297));
  INV_X1    g096(.A(new_n279), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n260), .A2(new_n264), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n284), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n283), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n294), .A2(new_n305), .A3(KEYINPUT70), .A4(new_n277), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT72), .A3(new_n283), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n295), .A2(new_n301), .B1(new_n305), .B2(new_n280), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n270), .A2(new_n282), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n316), .B2(new_n313), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n310), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G22gat), .ZN(new_n320));
  INV_X1    g119(.A(G228gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G141gat), .B(G148gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n328), .C1(new_n329), .C2(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G141gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n325), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(KEYINPUT2), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n330), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n343), .A3(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n324), .B1(new_n342), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n330), .A2(new_n338), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT29), .B1(new_n351), .B2(new_n352), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n354), .ZN(new_n364));
  INV_X1    g163(.A(new_n339), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n323), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n320), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  AOI211_X1 g168(.A(G22gat), .B(new_n367), .C1(new_n361), .C2(new_n362), .ZN(new_n370));
  OAI21_X1  g169(.A(G78gat), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n362), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT79), .B1(new_n355), .B2(new_n358), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G22gat), .ZN(new_n375));
  INV_X1    g174(.A(G78gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n363), .A2(new_n320), .A3(new_n368), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT31), .B(G50gat), .ZN(new_n380));
  INV_X1    g179(.A(G106gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(new_n378), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n341), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n243), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n215), .A2(new_n231), .A3(new_n242), .A4(new_n388), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n390), .A2(new_n353), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n353), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND4_X1  g196(.A1(new_n394), .A2(KEYINPUT74), .A3(KEYINPUT30), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n354), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n353), .A3(new_n391), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n401), .A4(new_n397), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n394), .A2(new_n397), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n330), .A2(new_n254), .A3(new_n258), .A4(new_n338), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT4), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n336), .B1(new_n337), .B2(new_n335), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n340), .A3(new_n259), .ZN(new_n417));
  NAND2_X1  g216(.A1(KEYINPUT77), .A2(KEYINPUT5), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n412), .A2(new_n413), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n330), .A4(new_n338), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n417), .A2(new_n420), .A3(new_n413), .A4(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n356), .A2(new_n259), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n431), .A2(new_n411), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n413), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n426), .A2(new_n430), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT81), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n419), .B2(new_n425), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n430), .A4(new_n437), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n430), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n435), .ZN(new_n444));
  INV_X1    g243(.A(new_n430), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n439), .A2(new_n442), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT82), .B(KEYINPUT35), .ZN(new_n448));
  NOR4_X1   g247(.A1(new_n386), .A2(new_n410), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n319), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n385), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n382), .B1(new_n371), .B2(new_n378), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n430), .A3(new_n435), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n436), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n430), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n438), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n405), .A3(new_n409), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n311), .A2(new_n314), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n310), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n310), .A2(new_n464), .A3(new_n315), .A4(new_n317), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n308), .A2(KEYINPUT72), .A3(new_n283), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT72), .B1(new_n308), .B2(new_n283), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n458), .B1(new_n384), .B2(new_n385), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n400), .A2(new_n401), .ZN(new_n472));
  INV_X1    g271(.A(new_n397), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n392), .B2(KEYINPUT80), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n400), .A2(new_n477), .A3(new_n401), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT38), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n397), .B1(new_n394), .B2(new_n475), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n473), .B1(new_n472), .B2(KEYINPUT37), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n394), .A2(new_n475), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT38), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n447), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n412), .A2(new_n417), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  INV_X1    g287(.A(new_n413), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n445), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n432), .A2(new_n413), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT39), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n487), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT39), .A3(new_n492), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(KEYINPUT40), .A3(new_n445), .A4(new_n490), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n495), .A2(new_n498), .A3(new_n454), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n410), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n471), .B1(new_n453), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n463), .B1(new_n470), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G197gat), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT11), .B(G169gat), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT12), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(KEYINPUT83), .A2(G36gat), .ZN(new_n511));
  OAI21_X1  g310(.A(G29gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT83), .B(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(G29gat), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  OR3_X1    g321(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT85), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n517), .A2(new_n521), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n513), .A3(new_n525), .A4(new_n516), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n520), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G1gat), .B2(new_n530), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G8gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n529), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT87), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT13), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n529), .A2(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT17), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT86), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT86), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n526), .A2(new_n528), .A3(new_n543), .A4(KEYINPUT17), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n534), .B1(new_n529), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n537), .B(new_n540), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n539), .B1(new_n548), .B2(KEYINPUT18), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n540), .B1(new_n545), .B2(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(new_n537), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n509), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n548), .A2(KEYINPUT18), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n508), .A4(new_n539), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n503), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(KEYINPUT92), .A2(G85gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G99gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT8), .B1(new_n578), .B2(new_n381), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n571), .A2(new_n577), .A3(new_n581), .A4(new_n579), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n529), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n529), .B2(new_n546), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n545), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n566), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n592), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n565), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n590), .A2(new_n566), .A3(new_n592), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n590), .A2(new_n592), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n601), .A2(new_n594), .A3(KEYINPUT93), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n590), .A2(KEYINPUT93), .A3(new_n592), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n564), .B(KEYINPUT91), .Z(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n599), .A2(new_n600), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G57gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT89), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT88), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n612), .A2(KEYINPUT88), .A3(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G71gat), .B(G78gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n611), .B(new_n617), .C1(new_n614), .C2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n534), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT90), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n584), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n619), .A3(new_n620), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n583), .A2(new_n584), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n645), .B2(KEYINPUT98), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n621), .A2(new_n641), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT97), .B(new_n654), .C1(new_n642), .C2(KEYINPUT10), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n585), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n619), .A3(new_n620), .A4(new_n639), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT10), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n656), .B1(new_n659), .B2(new_n653), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n643), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n651), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n653), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n645), .B1(new_n663), .B2(new_n644), .ZN(new_n664));
  INV_X1    g463(.A(new_n649), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n637), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n560), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n457), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT99), .B(G1gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1324gat));
  NAND3_X1  g471(.A1(new_n560), .A2(new_n410), .A3(new_n668), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT100), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(G8gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(new_n470), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n669), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n318), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n669), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n453), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  NOR3_X1   g486(.A1(new_n606), .A2(new_n636), .A3(new_n667), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n560), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n457), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n319), .A2(new_n449), .B1(new_n461), .B2(KEYINPUT35), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT102), .B1(new_n470), .B2(new_n502), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n501), .A2(new_n453), .ZN(new_n697));
  INV_X1    g496(.A(new_n471), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n469), .A4(new_n465), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n695), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n702), .B2(new_n606), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n602), .A2(new_n605), .ZN(new_n704));
  INV_X1    g503(.A(new_n600), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n598), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n503), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n636), .B(KEYINPUT101), .Z(new_n709));
  INV_X1    g508(.A(new_n559), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n710), .A3(new_n667), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n457), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(new_n410), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n514), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n689), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n514), .B1(new_n712), .B2(new_n715), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n470), .A3(new_n707), .A4(new_n711), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT47), .B1(new_n723), .B2(KEYINPUT103), .ZN(new_n724));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n689), .A2(new_n725), .A3(new_n319), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n724), .B(new_n727), .ZN(G1330gat));
  NAND4_X1  g527(.A1(new_n708), .A2(G50gat), .A3(new_n386), .A4(new_n711), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n560), .A2(new_n386), .A3(new_n688), .ZN(new_n730));
  INV_X1    g529(.A(G50gat), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(new_n731), .B1(KEYINPUT104), .B2(KEYINPUT48), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1331gat));
  INV_X1    g534(.A(new_n702), .ZN(new_n736));
  INV_X1    g535(.A(new_n667), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n637), .A2(new_n559), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n457), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n607), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n715), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n739), .A2(G71gat), .A3(new_n318), .ZN(new_n747));
  OAI21_X1  g546(.A(G71gat), .B1(new_n739), .B2(new_n681), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g549(.A1(new_n739), .A2(new_n453), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT105), .B(G78gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n574), .A2(new_n576), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n636), .A2(new_n559), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n737), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n708), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n754), .B1(new_n758), .B2(new_n457), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n702), .A2(new_n606), .A3(new_n756), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT106), .B(KEYINPUT51), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n737), .A2(new_n457), .A3(new_n754), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT107), .Z(new_n768));
  OAI21_X1  g567(.A(new_n759), .B1(new_n766), .B2(new_n768), .ZN(G1336gat));
  NOR3_X1   g568(.A1(new_n737), .A2(new_n715), .A3(G92gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n696), .A2(new_n701), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n606), .B1(new_n772), .B2(new_n463), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n773), .B2(new_n755), .ZN(new_n774));
  INV_X1    g573(.A(new_n771), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n702), .A2(new_n606), .A3(new_n756), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n770), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT109), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(new_n770), .C1(new_n774), .C2(new_n776), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n703), .A2(new_n410), .A3(new_n707), .A4(new_n757), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n765), .B2(new_n770), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n758), .B2(new_n681), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n318), .A2(new_n737), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n578), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n453), .A2(G106gat), .A3(new_n737), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT53), .B1(new_n765), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n703), .A2(new_n386), .A3(new_n707), .A4(new_n757), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n793), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n774), .A2(new_n776), .ZN(new_n799));
  INV_X1    g598(.A(new_n792), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n794), .A2(G106gat), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n803), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(new_n643), .C1(new_n659), .C2(new_n653), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n665), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n663), .B2(new_n644), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n806), .B(new_n809), .C1(new_n661), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n651), .A2(new_n661), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n661), .B2(new_n810), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n814), .A2(KEYINPUT55), .B1(new_n651), .B2(new_n661), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n661), .A2(new_n810), .ZN(new_n817));
  INV_X1    g616(.A(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n806), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n813), .A2(new_n559), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n550), .A2(new_n551), .B1(new_n535), .B2(new_n538), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n507), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n558), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n667), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n606), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n813), .A2(new_n820), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n706), .A2(new_n828), .A3(new_n824), .A4(new_n816), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n709), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n637), .A2(new_n559), .A3(new_n667), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n457), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n468), .A2(new_n386), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n715), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n246), .A3(new_n559), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n834), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n715), .A2(new_n691), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n386), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n319), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n710), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT112), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT112), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  AND4_X1   g645(.A1(G120gat), .A2(new_n839), .A3(new_n789), .A4(new_n841), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n837), .A2(new_n667), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n244), .ZN(G1341gat));
  NAND3_X1  g648(.A1(new_n837), .A2(new_n252), .A3(new_n636), .ZN(new_n850));
  OAI21_X1  g649(.A(G127gat), .B1(new_n842), .B2(new_n831), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1342gat));
  NOR3_X1   g651(.A1(new_n606), .A2(G134gat), .A3(new_n410), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n836), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n842), .B2(new_n606), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT113), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n470), .A2(new_n453), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n715), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n559), .A2(new_n331), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT118), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n470), .A2(new_n840), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT114), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n453), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n871));
  NAND2_X1  g670(.A1(new_n819), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n815), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n559), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n815), .B2(new_n872), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n825), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT117), .B(new_n825), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n606), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n636), .B1(new_n881), .B2(new_n829), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n870), .B1(new_n882), .B2(new_n833), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n709), .B1(new_n827), .B2(new_n829), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n386), .B1(new_n884), .B2(new_n833), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n869), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n710), .B(new_n868), .C1(new_n883), .C2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G141gat), .B1(new_n887), .B2(KEYINPUT120), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n868), .B1(new_n883), .B2(new_n886), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT120), .A3(new_n559), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n866), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n887), .A2(new_n331), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n892), .B2(new_n864), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(new_n861), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n333), .A3(new_n667), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n869), .B(new_n386), .C1(new_n882), .C2(new_n833), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n868), .A2(new_n737), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n333), .C1(new_n889), .C2(new_n667), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n896), .B1(new_n903), .B2(new_n904), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n895), .A2(new_n326), .A3(new_n636), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n889), .A2(new_n709), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n326), .ZN(G1346gat));
  NOR3_X1   g707(.A1(new_n606), .A2(G162gat), .A3(new_n410), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n835), .A2(new_n860), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n889), .A2(new_n706), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n327), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n410), .A2(new_n457), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n386), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n839), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n318), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n559), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G169gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n915), .A2(new_n468), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n202), .A3(new_n559), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1348gat));
  INV_X1    g723(.A(new_n920), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n203), .B1(new_n925), .B2(new_n737), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n839), .A2(G176gat), .A3(new_n789), .A4(new_n914), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT123), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n636), .A2(new_n228), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n225), .B1(new_n916), .B2(new_n709), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT60), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT60), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n229), .A3(new_n706), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n916), .A2(new_n706), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G190gat), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  NOR2_X1   g744(.A1(new_n470), .A2(new_n913), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n839), .A2(new_n386), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n948));
  XNOR2_X1  g747(.A(KEYINPUT125), .B(G197gat), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n839), .A2(new_n950), .A3(new_n386), .A4(new_n946), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n948), .A2(new_n559), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n946), .B(KEYINPUT126), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n900), .A2(new_n559), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n949), .ZN(G1352gat));
  NOR3_X1   g754(.A1(new_n947), .A2(G204gat), .A3(new_n737), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n900), .A2(new_n667), .A3(new_n953), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G204gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n900), .A2(new_n636), .A3(new_n953), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G211gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT63), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(new_n964), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(G211gat), .B1(new_n634), .B2(new_n635), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n951), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n963), .A2(new_n965), .A3(new_n968), .ZN(G1354gat));
  NAND4_X1  g768(.A1(new_n948), .A2(new_n346), .A3(new_n706), .A4(new_n951), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n900), .A2(new_n706), .A3(new_n953), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n346), .ZN(G1355gat));
endmodule


