//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT68), .A2(KEYINPUT23), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n213), .A2(G169gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n219), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n211), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT67), .B(G176gat), .Z(new_n226));
  AOI22_X1  g025(.A1(new_n226), .A2(new_n223), .B1(new_n217), .B2(new_n220), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n203), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n203), .A2(new_n228), .B1(new_n204), .B2(new_n205), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n207), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n207), .A2(new_n231), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n225), .B1(new_n235), .B2(KEYINPUT25), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n237), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n239));
  INV_X1    g038(.A(G120gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(G134gat), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n239), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G134gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(KEYINPUT72), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n249), .B2(new_n251), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n261));
  OAI221_X1 g060(.A(new_n216), .B1(KEYINPUT26), .B2(new_n220), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n205), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n264), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n236), .A2(new_n254), .A3(new_n258), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(new_n254), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n227), .B2(new_n234), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n211), .A2(new_n221), .A3(new_n224), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT64), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT33), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G43gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT73), .ZN(new_n282));
  XOR2_X1   g081(.A(G71gat), .B(G99gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n286));
  AOI221_X4 g085(.A(new_n286), .B1(KEYINPUT33), .B2(new_n284), .C1(new_n274), .C2(new_n276), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT34), .ZN(new_n289));
  INV_X1    g088(.A(new_n276), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n268), .A2(new_n273), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT34), .B1(new_n274), .B2(new_n276), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n285), .A2(new_n288), .A3(new_n293), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n295), .A3(new_n294), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n290), .B1(new_n268), .B2(new_n273), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n284), .B1(new_n299), .B2(KEYINPUT33), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n286), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n302), .B2(new_n287), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT86), .ZN(new_n307));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT2), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  OAI211_X1 g112(.A(KEYINPUT80), .B(new_n309), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(G148gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n315), .B1(new_n321), .B2(new_n309), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n329), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n323), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n330), .B(new_n332), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n316), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n315), .A3(new_n309), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n324), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n307), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT87), .ZN(new_n344));
  OR3_X1    g143(.A1(new_n337), .A2(new_n342), .A3(new_n306), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n307), .C1(new_n337), .C2(new_n342), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT88), .B1(new_n348), .B2(G22gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT31), .B(G50gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT89), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n349), .A2(KEYINPUT89), .A3(new_n353), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n348), .B(G22gat), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n357), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n349), .A2(KEYINPUT89), .A3(new_n353), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(new_n354), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n305), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n363));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n323), .B2(new_n336), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n339), .A2(new_n340), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n247), .A3(new_n253), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n258), .A2(new_n254), .A3(KEYINPUT4), .A4(new_n323), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n323), .B1(new_n256), .B2(new_n257), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n247), .A2(new_n367), .A3(new_n253), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n373), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n370), .B1(new_n366), .B2(new_n368), .ZN(new_n384));
  INV_X1    g183(.A(new_n379), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n384), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n258), .A2(new_n254), .A3(new_n376), .A4(new_n323), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n367), .B1(new_n247), .B2(new_n253), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n388), .A2(new_n389), .A3(new_n376), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT85), .B1(new_n375), .B2(KEYINPUT4), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n378), .A2(new_n383), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT84), .ZN(new_n395));
  XOR2_X1   g194(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n364), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT6), .B1(new_n393), .B2(new_n399), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n392), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n399), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n363), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n272), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n236), .A2(KEYINPUT79), .A3(new_n267), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n272), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n410), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n338), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n338), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n410), .B1(new_n413), .B2(new_n415), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n272), .B2(new_n324), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND3_X1  g224(.A1(new_n418), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n418), .A2(new_n422), .A3(KEYINPUT30), .A4(new_n425), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n202), .B1(new_n362), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n357), .B1(new_n355), .B2(new_n356), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n360), .A2(new_n359), .A3(new_n354), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n304), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(KEYINPUT96), .A3(new_n433), .A4(new_n409), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n302), .A2(new_n441), .A3(new_n287), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n298), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT74), .B1(new_n298), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n285), .A2(new_n288), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n404), .A2(new_n405), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n401), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(new_n408), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n440), .A2(new_n448), .A3(new_n452), .A4(new_n433), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n439), .B1(new_n453), .B2(KEYINPUT35), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n430), .A2(KEYINPUT37), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n338), .B1(new_n420), .B2(new_n421), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(KEYINPUT37), .C1(new_n460), .C2(new_n338), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(new_n426), .A3(new_n408), .A4(new_n407), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n429), .A2(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n458), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n440), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n392), .A2(new_n372), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT90), .B1(new_n469), .B2(new_n382), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471));
  AOI211_X1 g270(.A(new_n471), .B(new_n373), .C1(new_n392), .C2(new_n372), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT91), .A3(new_n399), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n389), .B1(new_n388), .B2(new_n376), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n375), .A2(KEYINPUT85), .A3(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n384), .B1(new_n478), .B2(new_n387), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n479), .B2(new_n373), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n258), .A2(new_n323), .A3(new_n254), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n376), .A2(new_n481), .B1(new_n476), .B2(new_n477), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT90), .B(new_n382), .C1(new_n482), .C2(new_n384), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT39), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n475), .B1(new_n484), .B2(new_n405), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n375), .A2(new_n373), .A3(new_n380), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n487), .B2(new_n486), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n474), .A2(new_n485), .A3(new_n490), .A4(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n400), .A2(new_n406), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n431), .A2(new_n432), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n428), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n485), .A3(new_n490), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT94), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  AND4_X1   g298(.A1(KEYINPUT94), .A2(new_n498), .A3(new_n491), .A4(new_n494), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n467), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n285), .A2(new_n288), .A3(KEYINPUT74), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n502), .A2(KEYINPUT76), .B1(new_n293), .B2(new_n296), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n293), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n504), .A2(KEYINPUT74), .B1(new_n285), .B2(new_n288), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT36), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n304), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n433), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n437), .B(new_n436), .C1(new_n510), .C2(new_n451), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n454), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(G1gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT16), .A3(new_n516), .ZN(new_n517));
  OAI221_X1 g316(.A(new_n517), .B1(KEYINPUT101), .B2(G8gat), .C1(new_n516), .C2(new_n515), .ZN(new_n518));
  NAND2_X1  g317(.A1(KEYINPUT101), .A2(G8gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G43gat), .B(G50gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n525), .B(KEYINPUT99), .Z(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NOR2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(new_n526), .A3(new_n528), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n531), .B2(new_n525), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT98), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n534), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n521), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n520), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n542), .A4(new_n544), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n543), .B(new_n520), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n542), .B(KEYINPUT13), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT97), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G169gat), .B(G197gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n547), .A2(new_n548), .A3(new_n551), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT102), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT102), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n514), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n576));
  AND2_X1   g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G127gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n520), .B1(KEYINPUT21), .B2(new_n575), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT103), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT104), .B(KEYINPUT7), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT105), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n598), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n599), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n600), .A2(KEYINPUT105), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n601), .A2(new_n603), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n608), .A2(new_n609), .A3(new_n604), .A4(new_n599), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n607), .B(new_n610), .C1(new_n539), .C2(new_n540), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT106), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n612), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n607), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n543), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n611), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n611), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n594), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n611), .A2(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n614), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n611), .A2(new_n615), .A3(new_n619), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n593), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n589), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n605), .A2(new_n606), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n605), .A2(new_n606), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n575), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n575), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n610), .A3(new_n607), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n636), .A2(KEYINPUT107), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n632), .A2(new_n634), .A3(new_n638), .A4(new_n635), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n629), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n632), .A2(new_n634), .ZN(new_n643));
  INV_X1    g442(.A(new_n629), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G120gat), .B(G148gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT108), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n642), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n568), .A2(new_n451), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g456(.A1(new_n628), .A2(new_n433), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n568), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n568), .A2(KEYINPUT109), .A3(new_n658), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(G8gat), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n661), .B2(new_n662), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n663), .B(new_n666), .C1(new_n667), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g467(.A1(new_n568), .A2(new_n655), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT36), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n444), .B2(new_n447), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n304), .A2(new_n507), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n506), .A2(KEYINPUT110), .A3(new_n508), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n304), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n669), .B2(new_n679), .ZN(G1326gat));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n358), .A2(new_n361), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n568), .A2(new_n683), .A3(new_n655), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n685), .A3(new_n681), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(G29gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n589), .A2(new_n627), .A3(new_n654), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n568), .A2(new_n692), .A3(new_n451), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n589), .B(KEYINPUT112), .ZN(new_n696));
  INV_X1    g495(.A(new_n654), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n562), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n514), .B2(new_n627), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n435), .A2(new_n439), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT94), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n496), .A2(new_n497), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n491), .A2(new_n494), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n498), .A2(KEYINPUT94), .A3(new_n491), .A4(new_n494), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n466), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n674), .A2(new_n511), .A3(new_n675), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n627), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n698), .B1(new_n699), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n452), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n695), .A2(new_n716), .ZN(G1328gat));
  NOR2_X1   g516(.A1(new_n433), .A2(G36gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n568), .A2(new_n693), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT46), .Z(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n715), .B2(new_n433), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n714), .B2(new_n676), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n702), .B1(new_n708), .B2(new_n512), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n304), .A2(G43gat), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n725), .A2(new_n566), .A3(new_n693), .A4(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT114), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI211_X1 g531(.A(KEYINPUT115), .B(KEYINPUT47), .C1(new_n727), .C2(KEYINPUT114), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n724), .A2(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n698), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n725), .B2(new_n711), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n676), .B(new_n735), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n730), .A2(new_n731), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT115), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(new_n729), .A3(new_n731), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n740), .A2(new_n742), .A3(new_n727), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(G1330gat));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  INV_X1    g545(.A(G50gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n714), .B2(new_n683), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n568), .A2(new_n747), .A3(new_n683), .A4(new_n693), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n683), .B(new_n735), .C1(new_n736), .C2(new_n738), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n749), .A3(KEYINPUT48), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1331gat));
  NOR3_X1   g554(.A1(new_n628), .A2(new_n562), .A3(new_n697), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n710), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n451), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g559(.A(new_n433), .B(KEYINPUT116), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n757), .B2(new_n677), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n304), .A2(G71gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n683), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n589), .A2(new_n562), .A3(new_n697), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n736), .B2(new_n738), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n452), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n589), .A2(new_n562), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n706), .A2(new_n707), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n709), .B1(new_n777), .B2(new_n467), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n711), .B(new_n776), .C1(new_n778), .C2(new_n454), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n711), .A4(new_n776), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n596), .A3(new_n451), .A4(new_n654), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n775), .A2(new_n784), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n774), .B2(new_n761), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n761), .A2(G92gat), .A3(new_n697), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n779), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n779), .B2(KEYINPUT117), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n510), .B(new_n773), .C1(new_n736), .C2(new_n738), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(new_n787), .B1(new_n793), .B2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n774), .B2(new_n677), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n697), .A2(new_n304), .A3(G99gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  OAI211_X1 g599(.A(new_n683), .B(new_n773), .C1(new_n736), .C2(new_n738), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n440), .A2(G106gat), .A3(new_n697), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT118), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n783), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n792), .A2(new_n804), .B1(new_n801), .B2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n636), .A2(KEYINPUT107), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n644), .A3(new_n640), .A4(new_n639), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n642), .A2(KEYINPUT119), .A3(KEYINPUT54), .A4(new_n811), .ZN(new_n815));
  INV_X1    g614(.A(new_n641), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n644), .B1(new_n816), .B2(new_n810), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n652), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n549), .A2(new_n550), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n542), .B1(new_n541), .B2(new_n544), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n557), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND4_X1   g624(.A1(new_n561), .A2(new_n622), .A3(new_n626), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n815), .A4(new_n819), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(new_n826), .A3(new_n653), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n827), .A2(new_n653), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT120), .A3(new_n822), .A4(new_n826), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n822), .A2(new_n562), .A3(new_n653), .A4(new_n827), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n654), .A2(new_n561), .A3(new_n825), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n711), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n696), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n562), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n655), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n761), .A2(new_n451), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n840), .A2(new_n362), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n567), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n452), .B1(new_n837), .B2(new_n839), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n440), .A2(new_n448), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n845), .A2(new_n847), .A3(new_n761), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n562), .A2(new_n242), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT121), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n851), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n848), .B2(new_n654), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n697), .A2(new_n240), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n842), .B2(new_n854), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n843), .B2(new_n696), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n848), .A2(new_n250), .A3(new_n589), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NOR2_X1   g657(.A1(new_n510), .A2(new_n627), .ZN(new_n859));
  XOR2_X1   g658(.A(KEYINPUT71), .B(G134gat), .Z(new_n860));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n847), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT56), .Z(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n843), .B2(new_n627), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n676), .A2(new_n841), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n837), .A2(new_n839), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n867), .B2(new_n683), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n683), .A2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n589), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n566), .A2(new_n822), .A3(new_n831), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n711), .B1(new_n871), .B2(new_n835), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(new_n833), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(new_n839), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n865), .B(G141gat), .C1(new_n875), .C2(new_n567), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n674), .A2(new_n683), .A3(new_n675), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT122), .Z(new_n878));
  NOR2_X1   g677(.A1(new_n567), .A2(G141gat), .ZN(new_n879));
  AND4_X1   g678(.A1(new_n761), .A2(new_n878), .A3(new_n845), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(KEYINPUT123), .B2(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n562), .B(new_n866), .C1(new_n868), .C2(new_n874), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n883), .A2(G141gat), .B1(new_n880), .B2(KEYINPUT123), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n865), .B2(new_n884), .ZN(G1344gat));
  AND2_X1   g684(.A1(new_n878), .A2(new_n845), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n761), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n887), .B2(new_n697), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n312), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n875), .A2(KEYINPUT59), .A3(new_n697), .ZN(new_n890));
  INV_X1    g689(.A(new_n828), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n870), .B1(new_n872), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n655), .A2(new_n567), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n683), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n840), .A2(new_n869), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n866), .A2(new_n654), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT59), .B(G148gat), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n889), .A2(new_n890), .A3(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n875), .B2(new_n696), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n870), .A2(G155gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n887), .B2(new_n902), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n875), .B2(new_n627), .ZN(new_n904));
  INV_X1    g703(.A(G162gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n905), .A3(new_n859), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n840), .A2(new_n362), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n451), .A2(new_n433), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n218), .A3(new_n567), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n867), .A2(new_n452), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n761), .B1(new_n912), .B2(KEYINPUT124), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n867), .A2(new_n914), .A3(new_n452), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n847), .A3(new_n562), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(new_n917), .B2(new_n218), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n910), .A2(new_n226), .A3(new_n697), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n847), .A3(new_n654), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n219), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n589), .A2(new_n263), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n913), .A2(new_n847), .A3(new_n915), .A4(new_n923), .ZN(new_n924));
  OR2_X1    g723(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n925));
  INV_X1    g724(.A(new_n696), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n867), .A2(new_n438), .A3(new_n926), .A4(new_n909), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n927), .A2(G183gat), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n924), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n711), .A3(new_n909), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(G190gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n933), .B2(G190gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n847), .A3(new_n915), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n711), .A2(new_n205), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  INV_X1    g738(.A(new_n877), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n916), .A2(new_n562), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n677), .A2(new_n909), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT126), .Z(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n897), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n567), .A2(new_n942), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n941), .A2(new_n942), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n913), .A2(new_n940), .A3(new_n915), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT127), .B(G204gat), .Z(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n697), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n949), .A2(KEYINPUT62), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n944), .B1(new_n895), .B2(new_n896), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(new_n697), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT62), .B1(new_n949), .B2(new_n953), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(G1353gat));
  NAND4_X1  g757(.A1(new_n916), .A2(new_n327), .A3(new_n589), .A4(new_n940), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n589), .B(new_n944), .C1(new_n895), .C2(new_n896), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n955), .B2(new_n627), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n711), .A2(new_n328), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n949), .B2(new_n965), .ZN(G1355gat));
endmodule


