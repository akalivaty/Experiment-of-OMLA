

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U552 ( .A1(n724), .A2(n723), .ZN(n731) );
  BUF_X1 U553 ( .A(n901), .Z(n518) );
  BUF_X1 U554 ( .A(n901), .Z(n519) );
  XNOR2_X1 U555 ( .A(n524), .B(n523), .ZN(n901) );
  NOR2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NAND2_X1 U557 ( .A1(n901), .A2(G137), .ZN(n553) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n625) );
  INV_X1 U559 ( .A(KEYINPUT68), .ZN(n554) );
  OR2_X1 U560 ( .A1(n728), .A2(n722), .ZN(n520) );
  NOR2_X1 U561 ( .A1(n719), .A2(n728), .ZN(n521) );
  XOR2_X1 U562 ( .A(KEYINPUT65), .B(n721), .Z(n522) );
  AND2_X1 U563 ( .A1(n645), .A2(n644), .ZN(n657) );
  INV_X1 U564 ( .A(KEYINPUT100), .ZN(n655) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n683) );
  INV_X1 U566 ( .A(KEYINPUT31), .ZN(n696) );
  BUF_X1 U567 ( .A(n659), .Z(n700) );
  NOR2_X1 U568 ( .A1(G1966), .A2(n728), .ZN(n712) );
  AND2_X1 U569 ( .A1(n720), .A2(n521), .ZN(n721) );
  NAND2_X1 U570 ( .A1(n520), .A2(n984), .ZN(n723) );
  NOR2_X1 U571 ( .A1(n733), .A2(n732), .ZN(n734) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U573 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n527), .ZN(n896) );
  XNOR2_X1 U575 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n752) );
  AND2_X1 U576 ( .A1(n560), .A2(n559), .ZN(G160) );
  INV_X1 U577 ( .A(G2105), .ZN(n527) );
  AND2_X1 U578 ( .A1(n527), .A2(G2104), .ZN(n900) );
  NAND2_X1 U579 ( .A1(G102), .A2(n900), .ZN(n526) );
  NAND2_X1 U580 ( .A1(G138), .A2(n519), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G126), .A2(n896), .ZN(n529) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U584 ( .A1(G114), .A2(n897), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n531), .A2(n530), .ZN(G164) );
  NOR2_X1 U587 ( .A1(G543), .A2(G651), .ZN(n794) );
  NAND2_X1 U588 ( .A1(n794), .A2(G89), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n587) );
  INV_X1 U591 ( .A(G651), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n587), .A2(n536), .ZN(n795) );
  NAND2_X1 U593 ( .A1(G76), .A2(n795), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n535), .B(KEYINPUT5), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(n536), .ZN(n538) );
  XNOR2_X1 U597 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n537) );
  XNOR2_X2 U598 ( .A(n538), .B(n537), .ZN(n790) );
  NAND2_X1 U599 ( .A1(G63), .A2(n790), .ZN(n541) );
  NOR2_X1 U600 ( .A1(n587), .A2(G651), .ZN(n539) );
  XOR2_X1 U601 ( .A(KEYINPUT67), .B(n539), .Z(n791) );
  NAND2_X1 U602 ( .A1(G51), .A2(n791), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G85), .A2(n794), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G72), .A2(n795), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G60), .A2(n790), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G47), .A2(n791), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U614 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U615 ( .A1(G113), .A2(n897), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n896), .A2(G125), .ZN(n556) );
  AND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G101), .A2(n900), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT23), .B(n558), .Z(n559) );
  NAND2_X1 U622 ( .A1(G61), .A2(n790), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G86), .A2(n794), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n795), .A2(G73), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT2), .B(n563), .Z(n564) );
  NOR2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n791), .A2(G48), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(G305) );
  NAND2_X1 U630 ( .A1(n791), .A2(G52), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT70), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G64), .A2(n790), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G90), .A2(n794), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G77), .A2(n795), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U639 ( .A1(n794), .A2(G88), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT82), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G75), .A2(n795), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT83), .B(n579), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G62), .A2(n790), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G50), .A2(n791), .ZN(n580) );
  AND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(G303) );
  NAND2_X1 U648 ( .A1(G49), .A2(n791), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n790), .A2(n586), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(G87), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(G288) );
  XOR2_X1 U654 ( .A(G1986), .B(KEYINPUT88), .Z(n590) );
  XNOR2_X1 U655 ( .A(G290), .B(n590), .ZN(n968) );
  NAND2_X1 U656 ( .A1(G105), .A2(n900), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n591), .B(KEYINPUT38), .ZN(n598) );
  NAND2_X1 U658 ( .A1(G141), .A2(n519), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G117), .A2(n897), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n896), .A2(G129), .ZN(n594) );
  XOR2_X1 U662 ( .A(KEYINPUT94), .B(n594), .Z(n595) );
  NOR2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n881) );
  NAND2_X1 U665 ( .A1(G1996), .A2(n881), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT95), .B(n599), .ZN(n610) );
  NAND2_X1 U667 ( .A1(G131), .A2(n518), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT92), .ZN(n607) );
  NAND2_X1 U669 ( .A1(G119), .A2(n896), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G107), .A2(n897), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G95), .A2(n900), .ZN(n603) );
  XNOR2_X1 U673 ( .A(KEYINPUT91), .B(n603), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n882) );
  NAND2_X1 U676 ( .A1(G1991), .A2(n882), .ZN(n608) );
  XNOR2_X1 U677 ( .A(KEYINPUT93), .B(n608), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n927) );
  NAND2_X1 U679 ( .A1(n968), .A2(n927), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G160), .A2(G40), .ZN(n611) );
  NOR2_X1 U681 ( .A1(n625), .A2(n611), .ZN(n748) );
  NAND2_X1 U682 ( .A1(n612), .A2(n748), .ZN(n624) );
  XNOR2_X1 U683 ( .A(G2067), .B(KEYINPUT37), .ZN(n745) );
  NAND2_X1 U684 ( .A1(G104), .A2(n900), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G140), .A2(n518), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U687 ( .A(KEYINPUT34), .B(n615), .ZN(n622) );
  XNOR2_X1 U688 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n897), .A2(G116), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n896), .A2(G128), .ZN(n616) );
  XOR2_X1 U691 ( .A(KEYINPUT89), .B(n616), .Z(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U693 ( .A(n620), .B(n619), .Z(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT36), .B(n623), .ZN(n893) );
  NOR2_X1 U696 ( .A1(n745), .A2(n893), .ZN(n929) );
  NAND2_X1 U697 ( .A1(n748), .A2(n929), .ZN(n742) );
  NAND2_X1 U698 ( .A1(n624), .A2(n742), .ZN(n735) );
  AND2_X1 U699 ( .A1(n625), .A2(G40), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G160), .A2(n626), .ZN(n627) );
  XNOR2_X2 U701 ( .A(n627), .B(KEYINPUT64), .ZN(n659) );
  NAND2_X1 U702 ( .A1(n659), .A2(G8), .ZN(n728) );
  NOR2_X1 U703 ( .A1(G1981), .A2(G305), .ZN(n628) );
  XOR2_X1 U704 ( .A(n628), .B(KEYINPUT24), .Z(n629) );
  NOR2_X1 U705 ( .A1(n728), .A2(n629), .ZN(n733) );
  INV_X1 U706 ( .A(G1996), .ZN(n947) );
  NOR2_X1 U707 ( .A1(n659), .A2(n947), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(n645) );
  AND2_X1 U710 ( .A1(n659), .A2(G1341), .ZN(n643) );
  XOR2_X1 U711 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n633) );
  NAND2_X1 U712 ( .A1(G56), .A2(n790), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n633), .B(n632), .ZN(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n794), .A2(G81), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT12), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G68), .A2(n795), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n791), .A2(G43), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n970) );
  NOR2_X1 U723 ( .A1(n643), .A2(n970), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G79), .A2(n795), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n646), .B(KEYINPUT76), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G92), .A2(n794), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G54), .A2(n791), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G66), .A2(n790), .ZN(n649) );
  XNOR2_X1 U730 ( .A(KEYINPUT75), .B(n649), .ZN(n650) );
  NOR2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(KEYINPUT15), .B(n654), .ZN(n983) );
  NOR2_X1 U734 ( .A1(n657), .A2(n983), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n657), .A2(n983), .ZN(n663) );
  INV_X1 U737 ( .A(n659), .ZN(n685) );
  AND2_X1 U738 ( .A1(n685), .A2(G2067), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(KEYINPUT99), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n700), .A2(G1348), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U744 ( .A1(G2072), .A2(n685), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT27), .ZN(n668) );
  AND2_X1 U746 ( .A1(n700), .A2(G1956), .ZN(n667) );
  NOR2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n677) );
  NAND2_X1 U748 ( .A1(G65), .A2(n790), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G53), .A2(n791), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G91), .A2(n794), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G78), .A2(n795), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n804) );
  NAND2_X1 U755 ( .A1(n677), .A2(n804), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n682) );
  NOR2_X1 U757 ( .A1(n677), .A2(n804), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT28), .B(KEYINPUT98), .ZN(n678) );
  XNOR2_X1 U759 ( .A(n678), .B(KEYINPUT97), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U762 ( .A(n684), .B(n683), .ZN(n689) );
  XNOR2_X1 U763 ( .A(KEYINPUT25), .B(G2078), .ZN(n946) );
  NAND2_X1 U764 ( .A1(n685), .A2(n946), .ZN(n687) );
  INV_X1 U765 ( .A(G1961), .ZN(n994) );
  NAND2_X1 U766 ( .A1(n700), .A2(n994), .ZN(n686) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n693), .A2(G171), .ZN(n688) );
  NAND2_X1 U769 ( .A1(n689), .A2(n688), .ZN(n699) );
  NOR2_X1 U770 ( .A1(n700), .A2(G2084), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n712), .A2(n708), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G8), .A2(n690), .ZN(n691) );
  XNOR2_X1 U773 ( .A(KEYINPUT30), .B(n691), .ZN(n692) );
  NOR2_X1 U774 ( .A1(G168), .A2(n692), .ZN(n695) );
  NOR2_X1 U775 ( .A1(G171), .A2(n693), .ZN(n694) );
  NOR2_X1 U776 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U777 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n710), .A2(G286), .ZN(n705) );
  NOR2_X1 U780 ( .A1(n700), .A2(G2090), .ZN(n702) );
  NOR2_X1 U781 ( .A1(G1971), .A2(n728), .ZN(n701) );
  NOR2_X1 U782 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U783 ( .A1(n703), .A2(G303), .ZN(n704) );
  NAND2_X1 U784 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U785 ( .A1(n706), .A2(G8), .ZN(n707) );
  XNOR2_X1 U786 ( .A(n707), .B(KEYINPUT32), .ZN(n716) );
  NAND2_X1 U787 ( .A1(G8), .A2(n708), .ZN(n709) );
  XNOR2_X1 U788 ( .A(KEYINPUT96), .B(n709), .ZN(n714) );
  INV_X1 U789 ( .A(n710), .ZN(n711) );
  NOR2_X1 U790 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U791 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U792 ( .A1(n716), .A2(n715), .ZN(n727) );
  NOR2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U794 ( .A1(G1971), .A2(G303), .ZN(n717) );
  NOR2_X1 U795 ( .A1(n971), .A2(n717), .ZN(n718) );
  NAND2_X1 U796 ( .A1(n727), .A2(n718), .ZN(n720) );
  NAND2_X1 U797 ( .A1(G1976), .A2(G288), .ZN(n972) );
  INV_X1 U798 ( .A(n972), .ZN(n719) );
  NOR2_X1 U799 ( .A1(KEYINPUT33), .A2(n522), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n971), .A2(KEYINPUT33), .ZN(n722) );
  XOR2_X1 U801 ( .A(G1981), .B(G305), .Z(n984) );
  NOR2_X1 U802 ( .A1(G2090), .A2(G303), .ZN(n725) );
  NAND2_X1 U803 ( .A1(G8), .A2(n725), .ZN(n726) );
  NAND2_X1 U804 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U807 ( .A(n736), .B(KEYINPUT101), .ZN(n751) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n881), .ZN(n922) );
  INV_X1 U809 ( .A(n927), .ZN(n739) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n882), .ZN(n918) );
  NOR2_X1 U812 ( .A1(n737), .A2(n918), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n922), .A2(n740), .ZN(n741) );
  XNOR2_X1 U815 ( .A(n741), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U817 ( .A(n744), .B(KEYINPUT102), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n745), .A2(n893), .ZN(n931) );
  NAND2_X1 U819 ( .A1(n746), .A2(n931), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U821 ( .A(KEYINPUT103), .B(n749), .Z(n750) );
  NAND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U823 ( .A(n753), .B(n752), .ZN(G329) );
  XOR2_X1 U824 ( .A(G2430), .B(G2443), .Z(n755) );
  XNOR2_X1 U825 ( .A(KEYINPUT105), .B(G2451), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n755), .B(n754), .ZN(n762) );
  XOR2_X1 U827 ( .A(G2435), .B(G2427), .Z(n757) );
  XNOR2_X1 U828 ( .A(G2446), .B(G2454), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U830 ( .A(n758), .B(G2438), .Z(n760) );
  XNOR2_X1 U831 ( .A(G1348), .B(G1341), .ZN(n759) );
  XNOR2_X1 U832 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n762), .B(n761), .ZN(n763) );
  AND2_X1 U834 ( .A1(n763), .A2(G14), .ZN(G401) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(n804), .ZN(G299) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n831) );
  NAND2_X1 U841 ( .A1(n831), .A2(G567), .ZN(n765) );
  XNOR2_X1 U842 ( .A(n765), .B(KEYINPUT71), .ZN(n766) );
  XNOR2_X1 U843 ( .A(KEYINPUT11), .B(n766), .ZN(G234) );
  XOR2_X1 U844 ( .A(G860), .B(KEYINPUT74), .Z(n773) );
  OR2_X1 U845 ( .A1(n773), .A2(n970), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  NOR2_X1 U847 ( .A1(n983), .A2(G868), .ZN(n767) );
  XNOR2_X1 U848 ( .A(n767), .B(KEYINPUT77), .ZN(n769) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n768) );
  NAND2_X1 U850 ( .A1(n769), .A2(n768), .ZN(G284) );
  INV_X1 U851 ( .A(G868), .ZN(n770) );
  NOR2_X1 U852 ( .A1(G286), .A2(n770), .ZN(n772) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n771) );
  NOR2_X1 U854 ( .A1(n772), .A2(n771), .ZN(G297) );
  NAND2_X1 U855 ( .A1(n773), .A2(G559), .ZN(n774) );
  NAND2_X1 U856 ( .A1(n774), .A2(n983), .ZN(n775) );
  XNOR2_X1 U857 ( .A(n775), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n970), .ZN(n778) );
  NAND2_X1 U859 ( .A1(n983), .A2(G868), .ZN(n776) );
  NOR2_X1 U860 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U862 ( .A1(n896), .A2(G123), .ZN(n780) );
  XNOR2_X1 U863 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n780), .B(n779), .ZN(n787) );
  NAND2_X1 U865 ( .A1(G99), .A2(n900), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G111), .A2(n897), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G135), .A2(n519), .ZN(n783) );
  XNOR2_X1 U869 ( .A(KEYINPUT79), .B(n783), .ZN(n784) );
  NOR2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n919) );
  XNOR2_X1 U872 ( .A(G2096), .B(n919), .ZN(n788) );
  NOR2_X1 U873 ( .A1(G2100), .A2(n788), .ZN(n789) );
  XOR2_X1 U874 ( .A(KEYINPUT80), .B(n789), .Z(G156) );
  NAND2_X1 U875 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U878 ( .A1(G93), .A2(n794), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G80), .A2(n795), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U881 ( .A1(n799), .A2(n798), .ZN(n811) );
  NAND2_X1 U882 ( .A1(n983), .A2(G559), .ZN(n814) );
  XNOR2_X1 U883 ( .A(n970), .B(n814), .ZN(n800) );
  NOR2_X1 U884 ( .A1(G860), .A2(n800), .ZN(n801) );
  XOR2_X1 U885 ( .A(KEYINPUT81), .B(n801), .Z(n802) );
  XNOR2_X1 U886 ( .A(n811), .B(n802), .ZN(G145) );
  INV_X1 U887 ( .A(G303), .ZN(G166) );
  NOR2_X1 U888 ( .A1(G868), .A2(n811), .ZN(n803) );
  XOR2_X1 U889 ( .A(n803), .B(KEYINPUT86), .Z(n817) );
  XNOR2_X1 U890 ( .A(n804), .B(G290), .ZN(n813) );
  XNOR2_X1 U891 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n806) );
  XNOR2_X1 U892 ( .A(G288), .B(KEYINPUT85), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G166), .B(n807), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(n970), .ZN(n809) );
  XOR2_X1 U896 ( .A(G305), .B(n809), .Z(n810) );
  XNOR2_X1 U897 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n862) );
  XNOR2_X1 U899 ( .A(n862), .B(n814), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G868), .A2(n815), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U906 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U908 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n823) );
  NAND2_X1 U909 ( .A1(G132), .A2(G82), .ZN(n822) );
  XNOR2_X1 U910 ( .A(n823), .B(n822), .ZN(n824) );
  NOR2_X1 U911 ( .A1(n824), .A2(G218), .ZN(n825) );
  NAND2_X1 U912 ( .A1(G96), .A2(n825), .ZN(n837) );
  NAND2_X1 U913 ( .A1(n837), .A2(G2106), .ZN(n829) );
  NAND2_X1 U914 ( .A1(G69), .A2(G120), .ZN(n826) );
  NOR2_X1 U915 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G108), .A2(n827), .ZN(n838) );
  NAND2_X1 U917 ( .A1(n838), .A2(G567), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n839) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n830) );
  NOR2_X1 U920 ( .A1(n839), .A2(n830), .ZN(n834) );
  NAND2_X1 U921 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n833) );
  XNOR2_X1 U926 ( .A(KEYINPUT106), .B(n833), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U928 ( .A(KEYINPUT107), .B(n836), .Z(G188) );
  INV_X1 U930 ( .A(G132), .ZN(G219) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n839), .ZN(G319) );
  XNOR2_X1 U938 ( .A(G1961), .B(KEYINPUT112), .ZN(n849) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1956), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U942 ( .A(G1981), .B(G1966), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2474), .B(KEYINPUT41), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U949 ( .A(G2096), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n861) );
  XOR2_X1 U952 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT110), .B(G2678), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2100), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(G227) );
  XOR2_X1 U962 ( .A(KEYINPUT117), .B(n862), .Z(n864) );
  XNOR2_X1 U963 ( .A(G171), .B(G286), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n983), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(G37), .A2(n866), .ZN(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT118), .B(n867), .ZN(G397) );
  NAND2_X1 U968 ( .A1(G124), .A2(n896), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G136), .A2(n518), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT113), .B(n869), .Z(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G100), .A2(n900), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G112), .A2(n897), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n919), .B(KEYINPUT116), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U980 ( .A(n878), .B(KEYINPUT114), .Z(n880) );
  XNOR2_X1 U981 ( .A(G164), .B(KEYINPUT115), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n885) );
  XNOR2_X1 U983 ( .A(G162), .B(n881), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n895) );
  NAND2_X1 U986 ( .A1(G103), .A2(n900), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G139), .A2(n519), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G127), .A2(n896), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G115), .A2(n897), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n933) );
  XNOR2_X1 U994 ( .A(n893), .B(n933), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n909) );
  NAND2_X1 U996 ( .A1(G130), .A2(n896), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G118), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U999 ( .A1(G106), .A2(n900), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n518), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT45), .B(n904), .Z(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(G160), .B(n907), .Z(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n913), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G397), .A2(G395), .ZN(n914) );
  XOR2_X1 U1012 ( .A(KEYINPUT119), .B(n914), .Z(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1016 ( .A(G160), .B(G2084), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n923), .B(KEYINPUT51), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n930), .B(KEYINPUT120), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n939) );
  XNOR2_X1 U1027 ( .A(G2072), .B(n933), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(G164), .B(G2078), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT121), .B(n936), .Z(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n937), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(n940), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT52), .ZN(n943) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT123), .B(n945), .Z(n1023) );
  XNOR2_X1 U1039 ( .A(G27), .B(n946), .ZN(n957) );
  XNOR2_X1 U1040 ( .A(G32), .B(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G28), .ZN(n955) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n953) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2072), .B(G33), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT124), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(KEYINPUT53), .ZN(n961) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n964), .ZN(n966) );
  INV_X1 U1057 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n967), .A2(G11), .ZN(n1021) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n982) );
  XNOR2_X1 U1063 ( .A(G1341), .B(n970), .ZN(n976) );
  INV_X1 U1064 ( .A(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(KEYINPUT126), .B(n974), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G299), .B(G1956), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G303), .B(G1971), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n991) );
  XOR2_X1 U1073 ( .A(G1348), .B(n983), .Z(n989) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(KEYINPUT125), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(KEYINPUT57), .B(n987), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1019) );
  INV_X1 U1081 ( .A(G16), .ZN(n1017) );
  XNOR2_X1 U1082 ( .A(G5), .B(n994), .ZN(n1012) );
  XNOR2_X1 U1083 ( .A(KEYINPUT59), .B(KEYINPUT127), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(G4), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1348), .B(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT60), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G21), .B(G1966), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

