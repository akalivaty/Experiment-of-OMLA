

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  XNOR2_X1 U321 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n443) );
  XNOR2_X1 U322 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U323 ( .A(n362), .B(n361), .ZN(n364) );
  XNOR2_X1 U324 ( .A(n419), .B(KEYINPUT120), .ZN(n420) );
  XNOR2_X1 U325 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U326 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U327 ( .A(n373), .B(n372), .Z(n569) );
  XNOR2_X1 U328 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U329 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(G71GAT), .B(KEYINPUT20), .Z(n294) );
  XOR2_X1 U331 ( .A(G99GAT), .B(KEYINPUT65), .Z(n290) );
  NAND2_X1 U332 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n292) );
  XNOR2_X1 U334 ( .A(G43GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n291), .B(G134GAT), .ZN(n399) );
  XNOR2_X1 U336 ( .A(n292), .B(n399), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n296) );
  XNOR2_X1 U338 ( .A(G15GAT), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(G127GAT), .ZN(n341) );
  XOR2_X1 U340 ( .A(n296), .B(n341), .Z(n302) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n298) );
  XNOR2_X1 U342 ( .A(KEYINPUT17), .B(G176GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(G169GAT), .B(n299), .Z(n325) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n300), .B(G120GAT), .ZN(n311) );
  XNOR2_X1 U347 ( .A(n325), .B(n311), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n532) );
  XOR2_X1 U349 ( .A(KEYINPUT4), .B(KEYINPUT86), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n323) );
  XOR2_X1 U352 ( .A(KEYINPUT78), .B(G85GAT), .Z(n306) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(G148GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT87), .B(G57GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(G127GAT), .B(G155GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(n310), .B(n309), .Z(n316) );
  XOR2_X1 U359 ( .A(G162GAT), .B(n311), .Z(n313) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(n314), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n317), .B(KEYINPUT1), .Z(n321) );
  XOR2_X1 U365 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n319) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(KEYINPUT82), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n430) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(n430), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n517) );
  XNOR2_X1 U371 ( .A(G8GAT), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n324), .B(G64GAT), .ZN(n340) );
  XOR2_X1 U373 ( .A(G36GAT), .B(G218GAT), .Z(n405) );
  XOR2_X1 U374 ( .A(n340), .B(n405), .Z(n327) );
  XOR2_X1 U375 ( .A(G197GAT), .B(KEYINPUT21), .Z(n427) );
  XNOR2_X1 U376 ( .A(n325), .B(n427), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U378 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n329) );
  NAND2_X1 U379 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U381 ( .A(n331), .B(n330), .Z(n336) );
  XOR2_X1 U382 ( .A(G92GAT), .B(G204GAT), .Z(n333) );
  XNOR2_X1 U383 ( .A(G183GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n334), .B(KEYINPUT89), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n473) );
  XOR2_X1 U387 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n338) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U390 ( .A(n339), .B(KEYINPUT80), .Z(n343) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U393 ( .A(n344), .B(KEYINPUT14), .Z(n346) );
  XOR2_X1 U394 ( .A(G22GAT), .B(G155GAT), .Z(n433) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(n433), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U397 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n348) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U400 ( .A(G57GAT), .B(n349), .Z(n385) );
  XNOR2_X1 U401 ( .A(n350), .B(n385), .ZN(n484) );
  INV_X1 U402 ( .A(n484), .ZN(n577) );
  XNOR2_X1 U403 ( .A(n577), .B(KEYINPUT110), .ZN(n565) );
  XOR2_X1 U404 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n391) );
  XOR2_X1 U405 ( .A(G1GAT), .B(G15GAT), .Z(n352) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G113GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n373) );
  XOR2_X1 U408 ( .A(G197GAT), .B(G141GAT), .Z(n354) );
  XNOR2_X1 U409 ( .A(G43GAT), .B(G22GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U411 ( .A(G36GAT), .B(G50GAT), .Z(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U413 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n358) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n360) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  INV_X1 U417 ( .A(KEYINPUT69), .ZN(n363) );
  NAND2_X1 U418 ( .A1(n364), .A2(n363), .ZN(n367) );
  INV_X1 U419 ( .A(n364), .ZN(n365) );
  NAND2_X1 U420 ( .A1(n365), .A2(KEYINPUT69), .ZN(n366) );
  NAND2_X1 U421 ( .A1(n367), .A2(n366), .ZN(n371) );
  XOR2_X1 U422 ( .A(G29GAT), .B(KEYINPUT8), .Z(n369) );
  XNOR2_X1 U423 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n400) );
  XNOR2_X1 U425 ( .A(n400), .B(KEYINPUT68), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U427 ( .A(G92GAT), .B(G85GAT), .Z(n375) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(G106GAT), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n403) );
  XOR2_X1 U430 ( .A(n403), .B(KEYINPUT76), .Z(n377) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n389) );
  XOR2_X1 U433 ( .A(KEYINPUT33), .B(G64GAT), .Z(n379) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G120GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U436 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U439 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U440 ( .A(G148GAT), .B(KEYINPUT75), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n384), .B(G204GAT), .ZN(n438) );
  XNOR2_X1 U442 ( .A(n438), .B(n385), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n573) );
  XNOR2_X1 U445 ( .A(KEYINPUT41), .B(n573), .ZN(n553) );
  AND2_X1 U446 ( .A1(n569), .A2(n553), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U448 ( .A1(n565), .A2(n392), .ZN(n410) );
  XOR2_X1 U449 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT9), .B(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n409) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n396) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n398) );
  INV_X1 U455 ( .A(KEYINPUT78), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n407) );
  XOR2_X1 U460 ( .A(G50GAT), .B(G162GAT), .Z(n429) );
  XOR2_X1 U461 ( .A(n429), .B(n405), .Z(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n559) );
  NAND2_X1 U464 ( .A1(n410), .A2(n559), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n411), .B(KEYINPUT47), .ZN(n417) );
  INV_X1 U466 ( .A(KEYINPUT36), .ZN(n412) );
  XNOR2_X1 U467 ( .A(KEYINPUT79), .B(n559), .ZN(n545) );
  XNOR2_X1 U468 ( .A(n412), .B(n545), .ZN(n584) );
  NOR2_X1 U469 ( .A1(n584), .A2(n484), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n413), .B(KEYINPUT45), .ZN(n414) );
  NAND2_X1 U471 ( .A1(n414), .A2(n573), .ZN(n415) );
  NOR2_X1 U472 ( .A1(n415), .A2(n569), .ZN(n416) );
  NOR2_X1 U473 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT48), .B(n418), .ZN(n530) );
  NOR2_X1 U475 ( .A1(n473), .A2(n530), .ZN(n421) );
  INV_X1 U476 ( .A(KEYINPUT54), .ZN(n419) );
  NOR2_X1 U477 ( .A1(n517), .A2(n422), .ZN(n568) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT85), .B(G78GAT), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n442) );
  XOR2_X1 U481 ( .A(KEYINPUT84), .B(G211GAT), .Z(n426) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(G106GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n436) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U490 ( .A(n437), .B(KEYINPUT23), .Z(n440) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT83), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n461) );
  NAND2_X1 U494 ( .A1(n568), .A2(n461), .ZN(n444) );
  NOR2_X1 U495 ( .A1(n532), .A2(n445), .ZN(n564) );
  NAND2_X1 U496 ( .A1(n564), .A2(n553), .ZN(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  NAND2_X1 U501 ( .A1(n564), .A2(n545), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n450) );
  XNOR2_X1 U503 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n472) );
  NAND2_X1 U504 ( .A1(n569), .A2(n573), .ZN(n487) );
  NOR2_X1 U505 ( .A1(n545), .A2(n484), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT16), .ZN(n470) );
  INV_X1 U507 ( .A(n532), .ZN(n523) );
  XNOR2_X1 U508 ( .A(n523), .B(KEYINPUT81), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n461), .B(KEYINPUT67), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT28), .ZN(n535) );
  XOR2_X1 U511 ( .A(n473), .B(KEYINPUT27), .Z(n463) );
  NAND2_X1 U512 ( .A1(n463), .A2(n517), .ZN(n529) );
  NOR2_X1 U513 ( .A1(n535), .A2(n529), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n456), .A2(n455), .ZN(n469) );
  INV_X1 U515 ( .A(n517), .ZN(n467) );
  NOR2_X1 U516 ( .A1(n532), .A2(n473), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT91), .B(n457), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n458), .A2(n461), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(KEYINPUT92), .Z(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n461), .A2(n523), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(n462), .ZN(n567) );
  NAND2_X1 U523 ( .A1(n567), .A2(n463), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n483) );
  NAND2_X1 U527 ( .A1(n470), .A2(n483), .ZN(n503) );
  NOR2_X1 U528 ( .A1(n487), .A2(n503), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n480), .A2(n517), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT93), .Z(n475) );
  INV_X1 U532 ( .A(n473), .ZN(n520) );
  NAND2_X1 U533 ( .A1(n480), .A2(n520), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT35), .B(KEYINPUT95), .Z(n477) );
  NAND2_X1 U536 ( .A1(n480), .A2(n523), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT94), .Z(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n480), .A2(n535), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n485), .A2(n584), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT37), .ZN(n516) );
  NOR2_X1 U547 ( .A1(n516), .A2(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT97), .B(n488), .Z(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n489), .ZN(n499) );
  NAND2_X1 U550 ( .A1(n499), .A2(n517), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n493) );
  NAND2_X1 U553 ( .A1(n499), .A2(n520), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n496) );
  NAND2_X1 U558 ( .A1(n499), .A2(n523), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n535), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT102), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  INV_X1 U564 ( .A(n569), .ZN(n502) );
  NAND2_X1 U565 ( .A1(n553), .A2(n502), .ZN(n515) );
  NOR2_X1 U566 ( .A1(n515), .A2(n503), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT103), .B(n504), .Z(n511) );
  NAND2_X1 U568 ( .A1(n517), .A2(n511), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n520), .A2(n511), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U575 ( .A1(n511), .A2(n523), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n535), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT107), .Z(n519) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n526), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  XOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n535), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT112), .B(n531), .Z(n551) );
  NOR2_X1 U597 ( .A1(n532), .A2(n551), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT113), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n569), .A2(n546), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U603 ( .A1(n546), .A2(n553), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT115), .Z(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U608 ( .A1(n546), .A2(n565), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  INV_X1 U615 ( .A(n567), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n569), .A2(n561), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n577), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n569), .A2(n564), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n583) );
  INV_X1 U635 ( .A(n583), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n575) );
  OR2_X1 U640 ( .A1(n583), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

