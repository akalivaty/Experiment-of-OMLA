//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT91), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT18), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G229gat), .A2(G233gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT87), .B(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G29gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n217), .C1(KEYINPUT15), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT88), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(G1gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n228), .A2(new_n231), .B1(KEYINPUT89), .B2(G8gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n227), .A3(new_n232), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT90), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n224), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n221), .B2(new_n222), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n239), .A2(KEYINPUT90), .B1(new_n234), .B2(new_n235), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n211), .B(new_n212), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n212), .B(KEYINPUT13), .Z(new_n242));
  INV_X1    g041(.A(new_n235), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n223), .B(KEYINPUT92), .C1(new_n243), .C2(new_n233), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n234), .A2(new_n235), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n223), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT92), .B1(new_n245), .B2(new_n223), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n209), .A2(new_n210), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(new_n212), .C1(new_n238), .C2(new_n240), .ZN(new_n251));
  INV_X1    g050(.A(new_n211), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI211_X1 g052(.A(KEYINPUT86), .B(new_n208), .C1(new_n249), .C2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n248), .A3(new_n241), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n207), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G231gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(G183gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G211gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT94), .B(KEYINPUT96), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G64gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT93), .A2(KEYINPUT9), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n270), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT20), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n245), .B1(new_n277), .B2(new_n276), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n279), .B(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n284), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n267), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n288), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n282), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n289), .A3(new_n266), .ZN(new_n296));
  NAND2_X1  g095(.A1(G99gat), .A2(G106gat), .ZN(new_n297));
  INV_X1    g096(.A(G85gat), .ZN(new_n298));
  INV_X1    g097(.A(G92gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(KEYINPUT8), .A2(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n298), .B2(new_n299), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT97), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G99gat), .B(G106gat), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n304), .B(KEYINPUT97), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n311), .A3(new_n237), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(new_n223), .ZN(new_n313));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT41), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n314), .B(KEYINPUT41), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G190gat), .B(G218gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G134gat), .B(G162gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  OR2_X1    g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n319), .A3(new_n323), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n309), .A2(new_n310), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n306), .A2(new_n307), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n275), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n276), .A2(new_n308), .A3(new_n311), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT10), .B(new_n275), .C1(new_n327), .C2(new_n328), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n329), .B2(new_n331), .ZN(new_n337));
  XOR2_X1   g136(.A(G120gat), .B(G148gat), .Z(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n335), .B(KEYINPUT100), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n332), .B2(new_n333), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n348), .B2(new_n337), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n292), .A2(new_n296), .A3(new_n326), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  OR2_X1    g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  INV_X1    g154(.A(G148gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G141gat), .ZN(new_n357));
  INV_X1    g156(.A(G141gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G148gat), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n355), .C1(new_n360), .C2(KEYINPUT2), .ZN(new_n361));
  OR2_X1    g160(.A1(KEYINPUT72), .A2(G162gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(KEYINPUT72), .A2(G162gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(G155gat), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT73), .A3(KEYINPUT2), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n357), .A2(new_n359), .B1(new_n354), .B2(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT73), .B1(new_n364), .B2(KEYINPUT2), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G113gat), .ZN(new_n371));
  INV_X1    g170(.A(G113gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G120gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G127gat), .B(G134gat), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  INV_X1    g182(.A(new_n380), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n375), .B2(new_n374), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n369), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n382), .B1(new_n389), .B2(KEYINPUT75), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  INV_X1    g190(.A(new_n363), .ZN(new_n392));
  NOR2_X1   g191(.A1(KEYINPUT72), .A2(G162gat), .ZN(new_n393));
  INV_X1    g192(.A(G155gat), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n365), .A3(new_n366), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n386), .A2(new_n387), .B1(new_n398), .B2(new_n361), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n353), .B1(new_n390), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT4), .B1(new_n369), .B2(new_n381), .ZN(new_n403));
  INV_X1    g202(.A(new_n381), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n398), .A4(new_n361), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n398), .A2(new_n409), .A3(new_n361), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n410), .A3(new_n388), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n407), .A2(new_n353), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT5), .B1(new_n402), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(new_n298), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n353), .A3(new_n411), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430));
  INV_X1    g229(.A(G190gat), .ZN(new_n431));
  AND2_X1   g230(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(G169gat), .A2(G176gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT26), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n436), .B(new_n431), .C1(new_n433), .C2(new_n432), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n438), .A2(new_n439), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT64), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n261), .A2(new_n431), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n449), .A2(new_n451), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(G169gat), .B2(G176gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458));
  INV_X1    g257(.A(G169gat), .ZN(new_n459));
  AND2_X1   g258(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT23), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n440), .B1(KEYINPUT23), .B2(new_n443), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n440), .A2(KEYINPUT23), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR3_X1    g266(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(new_n453), .A3(new_n448), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n458), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n430), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n447), .A4(new_n463), .ZN(new_n475));
  INV_X1    g274(.A(G226gat), .ZN(new_n476));
  INV_X1    g275(.A(G233gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(KEYINPUT29), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G218gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n263), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G204gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n203), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(G197gat), .A2(G204gat), .ZN(new_n488));
  OAI22_X1  g287(.A1(KEYINPUT22), .A2(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(G211gat), .B(G218gat), .Z(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n429), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  AOI211_X1 g294(.A(KEYINPUT70), .B(new_n495), .C1(new_n480), .C2(new_n482), .ZN(new_n496));
  INV_X1    g295(.A(new_n478), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n472), .B2(new_n475), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n447), .A3(new_n463), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n479), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n498), .A2(new_n501), .A3(new_n493), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n494), .A2(new_n496), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n428), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n483), .B2(new_n495), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n498), .A2(new_n501), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n493), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT38), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n483), .A2(new_n493), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n511));
  INV_X1    g310(.A(new_n498), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n495), .A3(new_n500), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n483), .A2(new_n429), .A3(new_n493), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n428), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n495), .B1(new_n480), .B2(new_n482), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n429), .A2(new_n517), .B1(new_n507), .B2(new_n495), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n511), .A4(new_n428), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n505), .A2(new_n509), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n522));
  INV_X1    g321(.A(new_n353), .ZN(new_n523));
  OAI22_X1  g322(.A1(new_n399), .A2(new_n400), .B1(new_n381), .B2(new_n369), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n389), .A2(KEYINPUT75), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n420), .B1(new_n526), .B2(new_n419), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n419), .A2(new_n420), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n417), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n424), .A2(new_n521), .A3(new_n522), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n419), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n528), .B1(new_n534), .B2(KEYINPUT5), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(new_n423), .A3(KEYINPUT6), .A4(new_n418), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n422), .A2(KEYINPUT76), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n504), .A3(new_n511), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n427), .A3(new_n509), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n519), .B1(new_n503), .B2(new_n428), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n514), .A2(new_n513), .ZN(new_n542));
  NOR4_X1   g341(.A1(new_n542), .A2(new_n494), .A3(KEYINPUT71), .A4(new_n427), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT85), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT37), .B1(new_n542), .B2(new_n494), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n505), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT38), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G50gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n369), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n493), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(new_n409), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n493), .B1(new_n410), .B2(new_n555), .ZN(new_n558));
  OAI211_X1 g357(.A(G228gat), .B(G233gat), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n561));
  OR3_X1    g360(.A1(new_n489), .A2(new_n561), .A3(new_n490), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n489), .B2(new_n490), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT79), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n489), .A2(new_n565), .A3(new_n490), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT3), .B1(new_n567), .B2(new_n555), .ZN(new_n568));
  INV_X1    g367(.A(G228gat), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n568), .A2(new_n554), .B1(new_n569), .B2(new_n477), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n559), .B(new_n560), .C1(new_n570), .C2(new_n558), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n558), .ZN(new_n573));
  OAI221_X1 g372(.A(new_n573), .B1(new_n569), .B2(new_n477), .C1(new_n554), .C2(new_n568), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n560), .B1(new_n574), .B2(new_n559), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT80), .B(new_n553), .C1(new_n572), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n559), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G22gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n553), .A2(KEYINPUT80), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n553), .A2(KEYINPUT80), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n571), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n427), .B1(new_n542), .B2(new_n494), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n515), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n516), .A2(new_n520), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n584), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n390), .A2(new_n353), .A3(new_n401), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT83), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT83), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n390), .A2(new_n591), .A3(new_n353), .A4(new_n401), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n353), .B1(new_n407), .B2(new_n411), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n590), .A2(KEYINPUT39), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n417), .B1(new_n596), .B2(KEYINPUT40), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(KEYINPUT40), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n530), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n595), .A2(new_n599), .B1(new_n596), .B2(KEYINPUT40), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n582), .B1(new_n588), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n549), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n576), .A2(new_n581), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n587), .B2(new_n538), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n481), .A2(new_n404), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n499), .A2(new_n381), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(G227gat), .A3(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(G227gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G15gat), .B(G43gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G99gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n616), .B(new_n617), .C1(new_n614), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n613), .A2(KEYINPUT32), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT34), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT34), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n613), .A2(KEYINPUT32), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n622), .A2(new_n627), .A3(new_n629), .A4(new_n624), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n631), .A2(KEYINPUT36), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT36), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT81), .B1(new_n609), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n586), .A2(new_n584), .ZN(new_n637));
  INV_X1    g436(.A(new_n585), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n538), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n582), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT81), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n633), .A2(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n607), .A2(new_n636), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n631), .A2(new_n632), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n582), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT35), .B1(new_n647), .B2(new_n639), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT35), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n649), .A3(new_n587), .A4(new_n538), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n259), .B(new_n352), .C1(new_n644), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n538), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g454(.A1(new_n652), .A2(new_n588), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n656), .B2(new_n226), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  MUX2_X1   g458(.A(KEYINPUT42), .B(new_n657), .S(new_n659), .Z(G1325gat));
  INV_X1    g459(.A(new_n645), .ZN(new_n661));
  AOI21_X1  g460(.A(G15gat), .B1(new_n652), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n635), .A2(G15gat), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n652), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n652), .A2(new_n582), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(G1327gat));
  AOI21_X1  g467(.A(new_n259), .B1(new_n644), .B2(new_n651), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n292), .A2(new_n296), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n351), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n326), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G29gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n653), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT45), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n326), .B1(new_n644), .B2(new_n651), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n609), .A2(new_n635), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n607), .A2(new_n679), .B1(new_n648), .B2(new_n650), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n326), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n324), .A2(KEYINPUT104), .A3(new_n325), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI22_X1  g485(.A1(new_n677), .A2(new_n678), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n254), .B2(new_n257), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n251), .A2(new_n252), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n241), .A2(new_n248), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n256), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n208), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n255), .A2(new_n256), .A3(new_n207), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(KEYINPUT102), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n671), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n687), .B2(new_n698), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n538), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n676), .B1(new_n705), .B2(new_n674), .ZN(G1328gat));
  INV_X1    g505(.A(new_n216), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n673), .A2(new_n707), .A3(new_n588), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n587), .B1(new_n701), .B2(new_n704), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n707), .ZN(G1329gat));
  NOR2_X1   g511(.A1(new_n645), .A2(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n669), .A2(new_n672), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT107), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n635), .B1(new_n700), .B2(new_n703), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(KEYINPUT47), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n687), .A2(new_n635), .A3(new_n698), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(KEYINPUT108), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(KEYINPUT108), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n717), .A2(KEYINPUT47), .B1(new_n721), .B2(new_n722), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n699), .B2(new_n608), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n608), .A2(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n673), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n582), .B1(new_n700), .B2(new_n703), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n728), .A2(G50gat), .B1(new_n673), .B2(new_n725), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g529(.A1(new_n292), .A2(new_n296), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n326), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n680), .A2(new_n732), .A3(new_n351), .A4(new_n696), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n653), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n588), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  AOI21_X1  g539(.A(G71gat), .B1(new_n733), .B2(new_n661), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n635), .A2(G71gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n733), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n582), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n351), .A3(new_n696), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n687), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(KEYINPUT109), .A3(new_n653), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G85gat), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n748), .B2(new_n653), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n607), .A2(new_n679), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n651), .ZN(new_n754));
  INV_X1    g553(.A(new_n326), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n697), .A2(new_n670), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n680), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n680), .B2(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n538), .A2(G85gat), .A3(new_n351), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n750), .A2(new_n751), .B1(new_n765), .B2(new_n767), .ZN(G1336gat));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n587), .A2(G92gat), .A3(new_n351), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n609), .B(new_n635), .C1(new_n549), .C2(new_n606), .ZN(new_n771));
  INV_X1    g570(.A(new_n651), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n757), .B(KEYINPUT51), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT110), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n757), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n752), .B1(new_n775), .B2(new_n759), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n769), .B(new_n770), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n643), .A2(new_n636), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n604), .A2(new_n603), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n601), .B2(new_n600), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n608), .B1(new_n780), .B2(new_n587), .ZN(new_n781));
  INV_X1    g580(.A(new_n548), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n424), .A2(new_n521), .A3(new_n532), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(KEYINPUT85), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n784), .B2(new_n533), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n651), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n678), .B1(new_n786), .B2(new_n755), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n680), .A2(new_n686), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n588), .B(new_n747), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n777), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n769), .B1(new_n764), .B2(new_n770), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n762), .A2(new_n773), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n789), .A2(G92gat), .B1(new_n794), .B2(new_n770), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n792), .A2(new_n793), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI221_X1 g597(.A(KEYINPUT113), .B1(new_n791), .B2(new_n795), .C1(new_n792), .C2(new_n793), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1337gat));
  NAND2_X1  g599(.A1(new_n748), .A2(new_n635), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G99gat), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n645), .A2(G99gat), .A3(new_n351), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n765), .B2(new_n803), .ZN(G1338gat));
  NAND2_X1  g603(.A1(new_n748), .A2(new_n582), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n608), .A2(G106gat), .A3(new_n351), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n765), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(KEYINPUT114), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n805), .A2(G106gat), .B1(new_n794), .B2(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n808), .A2(new_n810), .B1(new_n812), .B2(new_n807), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n332), .A2(new_n333), .A3(new_n347), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n336), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n342), .B1(new_n348), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n818), .A2(new_n819), .B1(new_n336), .B2(new_n344), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n689), .B2(new_n695), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n246), .A2(new_n247), .A3(new_n242), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n238), .A2(new_n212), .A3(new_n240), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n206), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n249), .A2(new_n253), .A3(new_n207), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n827), .A2(new_n350), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n684), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n822), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n683), .A3(new_n682), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n731), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n352), .A2(new_n696), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n588), .A2(new_n538), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n838), .A2(new_n647), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n372), .A3(new_n696), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n258), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(new_n372), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n350), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n731), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G127gat), .ZN(G1342gat));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(new_n755), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(G134gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n852), .B2(KEYINPUT56), .ZN(new_n853));
  OR4_X1    g652(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT56), .A4(G134gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(G134gat), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n635), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n838), .B2(new_n608), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n332), .A2(new_n333), .A3(new_n347), .ZN(new_n863));
  INV_X1    g662(.A(new_n335), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n332), .B2(new_n333), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n865), .A3(new_n816), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n334), .A2(new_n816), .A3(new_n346), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n343), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n819), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n345), .A4(new_n821), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n693), .A3(new_n694), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n820), .B2(new_n821), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n830), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n326), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n731), .B1(new_n875), .B2(new_n835), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT57), .B(new_n582), .C1(new_n876), .C2(new_n837), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n358), .B1(new_n878), .B2(new_n258), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n836), .A2(new_n837), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n582), .A3(new_n858), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n258), .A2(new_n358), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  INV_X1    g686(.A(new_n885), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n879), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n358), .B1(new_n878), .B2(new_n696), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT58), .B1(new_n890), .B2(new_n884), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n889), .A3(new_n891), .ZN(G1344gat));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n882), .B2(new_n351), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n356), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n582), .B(new_n860), .C1(new_n836), .C2(new_n837), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n326), .A2(new_n822), .A3(new_n833), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n874), .B2(new_n326), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n898), .A2(new_n731), .B1(new_n258), .B2(new_n352), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n582), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n350), .A3(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT59), .B(G148gat), .C1(new_n901), .C2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n878), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n351), .A2(KEYINPUT59), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n894), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(G1345gat));
  INV_X1    g707(.A(new_n882), .ZN(new_n909));
  AOI21_X1  g708(.A(G155gat), .B1(new_n909), .B2(new_n731), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n670), .A2(new_n394), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n878), .B2(new_n911), .ZN(G1346gat));
  NAND2_X1  g711(.A1(new_n362), .A2(new_n363), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n913), .A3(new_n755), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n906), .A2(new_n684), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n913), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n653), .A2(new_n587), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n646), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n838), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n459), .A3(new_n696), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT121), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n258), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n459), .B2(new_n923), .ZN(G1348gat));
  NAND2_X1  g723(.A1(new_n919), .A2(new_n350), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G176gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n460), .A2(new_n461), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n925), .ZN(G1349gat));
  NAND2_X1  g727(.A1(new_n919), .A2(new_n731), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G183gat), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n432), .A2(new_n433), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n929), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g732(.A(new_n431), .B1(new_n919), .B2(new_n755), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT61), .Z(new_n935));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n431), .A3(new_n683), .A4(new_n682), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n642), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n897), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n731), .B1(new_n875), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n352), .A2(new_n258), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n582), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n940), .B1(new_n946), .B2(new_n895), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n259), .ZN(new_n949));
  INV_X1    g748(.A(new_n938), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n881), .A2(new_n582), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n203), .A3(new_n696), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n953), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n350), .A2(new_n486), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(KEYINPUT62), .C1(new_n951), .C2(new_n955), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n958), .A2(new_n960), .B1(new_n957), .B2(new_n956), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT124), .B1(new_n947), .B2(new_n350), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT124), .A3(new_n350), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(G1353gat));
  AOI21_X1  g764(.A(new_n263), .B1(new_n947), .B2(new_n731), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n966), .B2(KEYINPUT63), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n731), .B(new_n939), .C1(new_n896), .C2(new_n900), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n971), .A3(KEYINPUT63), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n670), .B(new_n940), .C1(new_n946), .C2(new_n895), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n973), .B(new_n974), .C1(new_n975), .C2(new_n263), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n967), .A2(new_n970), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n952), .A2(new_n263), .A3(new_n731), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(new_n484), .B1(new_n951), .B2(new_n684), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n755), .A2(G218gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n948), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT127), .Z(G1355gat));
endmodule


