

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725;

  NOR2_X1 U368 ( .A1(G953), .A2(G237), .ZN(n493) );
  INV_X1 U369 ( .A(n651), .ZN(n581) );
  INV_X1 U370 ( .A(G953), .ZN(n712) );
  XNOR2_X2 U371 ( .A(n535), .B(n517), .ZN(n645) );
  XNOR2_X2 U372 ( .A(n445), .B(n444), .ZN(n535) );
  AND2_X1 U373 ( .A1(n384), .A2(n381), .ZN(n380) );
  XNOR2_X1 U374 ( .A(n468), .B(n369), .ZN(n700) );
  INV_X1 U375 ( .A(G107), .ZN(n417) );
  INV_X1 U376 ( .A(G116), .ZN(n374) );
  INV_X1 U377 ( .A(G122), .ZN(n370) );
  XNOR2_X1 U378 ( .A(n404), .B(n403), .ZN(n720) );
  XNOR2_X1 U379 ( .A(n583), .B(n430), .ZN(n666) );
  NAND2_X1 U380 ( .A1(n380), .A2(n377), .ZN(n543) );
  XNOR2_X1 U381 ( .A(n461), .B(n460), .ZN(n647) );
  XNOR2_X1 U382 ( .A(n701), .B(n467), .ZN(n442) );
  XNOR2_X1 U383 ( .A(n373), .B(n372), .ZN(n468) );
  XNOR2_X1 U384 ( .A(n433), .B(G110), .ZN(n701) );
  XNOR2_X1 U385 ( .A(n371), .B(n370), .ZN(n369) );
  XNOR2_X1 U386 ( .A(n374), .B(G113), .ZN(n373) );
  XNOR2_X1 U387 ( .A(n411), .B(G143), .ZN(n512) );
  XNOR2_X1 U388 ( .A(n417), .B(G104), .ZN(n433) );
  XNOR2_X1 U389 ( .A(G119), .B(KEYINPUT3), .ZN(n372) );
  XNOR2_X1 U390 ( .A(KEYINPUT16), .B(KEYINPUT74), .ZN(n371) );
  AND2_X2 U391 ( .A1(n395), .A2(n674), .ZN(n347) );
  XNOR2_X1 U392 ( .A(n512), .B(n410), .ZN(n438) );
  NOR2_X2 U393 ( .A1(n697), .A2(n446), .ZN(n394) );
  AND2_X1 U394 ( .A1(n386), .A2(KEYINPUT89), .ZN(n385) );
  NAND2_X1 U395 ( .A1(n635), .A2(n383), .ZN(n382) );
  NAND2_X1 U396 ( .A1(n349), .A2(n592), .ZN(n390) );
  INV_X1 U397 ( .A(n711), .ZN(n393) );
  INV_X1 U398 ( .A(KEYINPUT89), .ZN(n383) );
  NOR2_X1 U399 ( .A1(n564), .A2(n485), .ZN(n486) );
  NAND2_X1 U400 ( .A1(n388), .A2(n446), .ZN(n387) );
  INV_X1 U401 ( .A(n349), .ZN(n388) );
  OR2_X1 U402 ( .A1(n596), .A2(G902), .ZN(n409) );
  XNOR2_X1 U403 ( .A(n413), .B(n412), .ZN(n551) );
  XNOR2_X1 U404 ( .A(n526), .B(KEYINPUT72), .ZN(n412) );
  NOR2_X1 U405 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U406 ( .A(n720), .ZN(n402) );
  XNOR2_X1 U407 ( .A(n397), .B(n396), .ZN(n429) );
  XNOR2_X1 U408 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n397) );
  NAND2_X1 U409 ( .A1(n712), .A2(G224), .ZN(n396) );
  XNOR2_X1 U410 ( .A(n406), .B(G125), .ZN(n456) );
  INV_X1 U411 ( .A(G146), .ZN(n406) );
  INV_X1 U412 ( .A(KEYINPUT4), .ZN(n410) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n588) );
  INV_X1 U414 ( .A(KEYINPUT44), .ZN(n357) );
  NAND2_X1 U415 ( .A1(n400), .A2(n725), .ZN(n358) );
  AND2_X1 U416 ( .A1(n402), .A2(n618), .ZN(n400) );
  NOR2_X1 U417 ( .A1(n549), .A2(n550), .ZN(n419) );
  NOR2_X1 U418 ( .A1(n529), .A2(n541), .ZN(n530) );
  AND2_X2 U419 ( .A1(n395), .A2(n674), .ZN(n688) );
  NOR2_X1 U420 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U421 ( .A(KEYINPUT36), .ZN(n362) );
  NOR2_X1 U422 ( .A1(n521), .A2(n575), .ZN(n554) );
  NAND2_X1 U423 ( .A1(n489), .A2(n568), .ZN(n415) );
  NOR2_X1 U424 ( .A1(n488), .A2(n487), .ZN(n489) );
  INV_X1 U425 ( .A(n519), .ZN(n487) );
  INV_X1 U426 ( .A(KEYINPUT105), .ZN(n360) );
  INV_X1 U427 ( .A(n529), .ZN(n542) );
  NOR2_X1 U428 ( .A1(n535), .A2(n644), .ZN(n568) );
  XNOR2_X1 U429 ( .A(n559), .B(n398), .ZN(n636) );
  INV_X1 U430 ( .A(KEYINPUT38), .ZN(n398) );
  XNOR2_X1 U431 ( .A(KEYINPUT69), .B(G137), .ZN(n436) );
  XOR2_X1 U432 ( .A(G131), .B(G134), .Z(n437) );
  XOR2_X1 U433 ( .A(G146), .B(KEYINPUT97), .Z(n465) );
  XOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n491) );
  XNOR2_X1 U435 ( .A(G113), .B(G104), .ZN(n490) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n495) );
  XNOR2_X1 U437 ( .A(G143), .B(G131), .ZN(n497) );
  XOR2_X1 U438 ( .A(G146), .B(G140), .Z(n440) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n479) );
  XOR2_X1 U440 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n480) );
  AND2_X1 U441 ( .A1(n636), .A2(n635), .ZN(n634) );
  INV_X1 U442 ( .A(n636), .ZN(n414) );
  INV_X1 U443 ( .A(n382), .ZN(n375) );
  NAND2_X1 U444 ( .A1(n651), .A2(n635), .ZN(n478) );
  NOR2_X1 U445 ( .A1(n647), .A2(n520), .ZN(n533) );
  XNOR2_X1 U446 ( .A(n456), .B(n405), .ZN(n708) );
  XNOR2_X1 U447 ( .A(G140), .B(KEYINPUT10), .ZN(n405) );
  XNOR2_X1 U448 ( .A(G137), .B(G110), .ZN(n451) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n452) );
  XNOR2_X1 U450 ( .A(G119), .B(G128), .ZN(n454) );
  XOR2_X1 U451 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n505) );
  XNOR2_X1 U452 ( .A(G116), .B(G134), .ZN(n502) );
  XOR2_X1 U453 ( .A(G122), .B(G107), .Z(n503) );
  XNOR2_X1 U454 ( .A(n700), .B(n427), .ZN(n426) );
  XNOR2_X1 U455 ( .A(n429), .B(n456), .ZN(n427) );
  INV_X1 U456 ( .A(KEYINPUT45), .ZN(n420) );
  NAND2_X1 U457 ( .A1(n418), .A2(n351), .ZN(n711) );
  XNOR2_X1 U458 ( .A(n419), .B(KEYINPUT48), .ZN(n418) );
  INV_X1 U459 ( .A(n632), .ZN(n560) );
  XNOR2_X1 U460 ( .A(n543), .B(KEYINPUT19), .ZN(n566) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n529) );
  XNOR2_X1 U462 ( .A(n501), .B(G475), .ZN(n407) );
  OR2_X1 U463 ( .A1(n606), .A2(G902), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n528), .B(KEYINPUT40), .ZN(n723) );
  NOR2_X1 U465 ( .A1(n645), .A2(n523), .ZN(n630) );
  XNOR2_X1 U466 ( .A(n522), .B(n361), .ZN(n523) );
  XNOR2_X1 U467 ( .A(n362), .B(KEYINPUT109), .ZN(n361) );
  XNOR2_X1 U468 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n403) );
  AND2_X1 U469 ( .A1(n578), .A2(n577), .ZN(n404) );
  INV_X1 U470 ( .A(n654), .ZN(n367) );
  INV_X1 U471 ( .A(n415), .ZN(n525) );
  INV_X1 U472 ( .A(n647), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n603), .B(n356), .ZN(n604) );
  XNOR2_X1 U474 ( .A(n365), .B(n355), .ZN(n689) );
  NAND2_X1 U475 ( .A1(n347), .A2(G469), .ZN(n365) );
  INV_X1 U476 ( .A(KEYINPUT56), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n425), .B(n353), .ZN(n424) );
  AND2_X1 U478 ( .A1(n581), .A2(n401), .ZN(n348) );
  XOR2_X1 U479 ( .A(n435), .B(n434), .Z(n349) );
  AND2_X1 U480 ( .A1(n570), .A2(n633), .ZN(n350) );
  AND2_X1 U481 ( .A1(n724), .A2(n560), .ZN(n351) );
  NOR2_X1 U482 ( .A1(n612), .A2(n350), .ZN(n352) );
  XOR2_X1 U483 ( .A(n682), .B(n681), .Z(n353) );
  XNOR2_X1 U484 ( .A(KEYINPUT35), .B(KEYINPUT78), .ZN(n354) );
  XOR2_X1 U485 ( .A(n687), .B(n686), .Z(n355) );
  XOR2_X1 U486 ( .A(n602), .B(KEYINPUT122), .Z(n356) );
  NOR2_X1 U487 ( .A1(G952), .A2(n712), .ZN(n693) );
  INV_X1 U488 ( .A(n693), .ZN(n423) );
  NAND2_X1 U489 ( .A1(n359), .A2(n348), .ZN(n618) );
  XNOR2_X1 U490 ( .A(n589), .B(n360), .ZN(n359) );
  NAND2_X1 U491 ( .A1(n688), .A2(G475), .ZN(n608) );
  NAND2_X1 U492 ( .A1(n363), .A2(n524), .ZN(n550) );
  XNOR2_X1 U493 ( .A(n630), .B(KEYINPUT87), .ZN(n363) );
  NAND2_X1 U494 ( .A1(n595), .A2(KEYINPUT2), .ZN(n674) );
  NAND2_X1 U495 ( .A1(n482), .A2(G902), .ZN(n562) );
  XNOR2_X1 U496 ( .A(n481), .B(KEYINPUT75), .ZN(n482) );
  XNOR2_X1 U497 ( .A(n364), .B(n422), .ZN(G51) );
  NAND2_X1 U498 ( .A1(n424), .A2(n423), .ZN(n364) );
  XOR2_X2 U499 ( .A(KEYINPUT95), .B(n472), .Z(n709) );
  NAND2_X1 U500 ( .A1(n392), .A2(n594), .ZN(n395) );
  NAND2_X1 U501 ( .A1(n394), .A2(n393), .ZN(n392) );
  AND2_X2 U502 ( .A1(n587), .A2(n586), .ZN(n399) );
  XNOR2_X1 U503 ( .A(n366), .B(n611), .ZN(G60) );
  NOR2_X2 U504 ( .A1(n609), .A2(n693), .ZN(n366) );
  AND2_X1 U505 ( .A1(n572), .A2(n367), .ZN(n569) );
  AND2_X1 U506 ( .A1(n572), .A2(n581), .ZN(n567) );
  NAND2_X1 U507 ( .A1(n368), .A2(n572), .ZN(n585) );
  XNOR2_X2 U508 ( .A(n416), .B(KEYINPUT0), .ZN(n572) );
  INV_X1 U509 ( .A(n666), .ZN(n368) );
  INV_X1 U510 ( .A(n376), .ZN(n389) );
  NAND2_X1 U511 ( .A1(n376), .A2(n375), .ZN(n381) );
  NAND2_X1 U512 ( .A1(n391), .A2(n390), .ZN(n376) );
  NAND2_X1 U513 ( .A1(n389), .A2(n386), .ZN(n559) );
  NOR2_X1 U514 ( .A1(n635), .A2(n383), .ZN(n378) );
  NOR2_X1 U515 ( .A1(n386), .A2(n382), .ZN(n379) );
  NAND2_X1 U516 ( .A1(n385), .A2(n389), .ZN(n384) );
  OR2_X1 U517 ( .A1(n680), .A2(n387), .ZN(n386) );
  NAND2_X1 U518 ( .A1(n680), .A2(n349), .ZN(n391) );
  NOR2_X1 U519 ( .A1(n697), .A2(n711), .ZN(n595) );
  XNOR2_X2 U520 ( .A(n399), .B(n354), .ZN(n725) );
  NOR2_X1 U521 ( .A1(n580), .A2(n576), .ZN(n578) );
  XNOR2_X2 U522 ( .A(n409), .B(n475), .ZN(n651) );
  XNOR2_X2 U523 ( .A(G128), .B(KEYINPUT80), .ZN(n411) );
  NOR2_X2 U524 ( .A1(n566), .A2(n565), .ZN(n416) );
  XNOR2_X2 U525 ( .A(n421), .B(n420), .ZN(n697) );
  NAND2_X1 U526 ( .A1(n588), .A2(n352), .ZN(n421) );
  NAND2_X1 U527 ( .A1(n347), .A2(G210), .ZN(n425) );
  XNOR2_X1 U528 ( .A(n428), .B(n426), .ZN(n680) );
  XNOR2_X1 U529 ( .A(n438), .B(n442), .ZN(n428) );
  XNOR2_X1 U530 ( .A(n598), .B(n597), .ZN(n599) );
  NOR2_X2 U531 ( .A1(n599), .A2(n693), .ZN(n601) );
  XNOR2_X1 U532 ( .A(n605), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U533 ( .A1(n604), .A2(n423), .ZN(n605) );
  NAND2_X1 U534 ( .A1(n688), .A2(G472), .ZN(n598) );
  INV_X1 U535 ( .A(n535), .ZN(n536) );
  XNOR2_X1 U536 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n430) );
  AND2_X1 U537 ( .A1(G221), .A2(n508), .ZN(n431) );
  XOR2_X1 U538 ( .A(n437), .B(n436), .Z(n432) );
  XNOR2_X1 U539 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U540 ( .A(G472), .ZN(n473) );
  XOR2_X1 U541 ( .A(n471), .B(n472), .Z(n596) );
  INV_X1 U542 ( .A(KEYINPUT34), .ZN(n584) );
  XNOR2_X1 U543 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U544 ( .A(n596), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U545 ( .A(n459), .B(n458), .ZN(n691) );
  INV_X1 U546 ( .A(KEYINPUT63), .ZN(n600) );
  XNOR2_X1 U547 ( .A(n601), .B(n600), .ZN(G57) );
  XNOR2_X1 U548 ( .A(G902), .B(KEYINPUT15), .ZN(n446) );
  INV_X1 U549 ( .A(n446), .ZN(n592) );
  XOR2_X1 U550 ( .A(KEYINPUT68), .B(G101), .Z(n467) );
  OR2_X1 U551 ( .A1(G237), .A2(G902), .ZN(n476) );
  NAND2_X1 U552 ( .A1(G210), .A2(n476), .ZN(n435) );
  XOR2_X1 U553 ( .A(KEYINPUT81), .B(KEYINPUT90), .Z(n434) );
  INV_X1 U554 ( .A(n559), .ZN(n516) );
  XNOR2_X1 U555 ( .A(n438), .B(n432), .ZN(n472) );
  NAND2_X1 U556 ( .A1(G227), .A2(n712), .ZN(n439) );
  XNOR2_X1 U557 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U558 ( .A(n709), .B(n443), .ZN(n685) );
  NOR2_X1 U559 ( .A1(G902), .A2(n685), .ZN(n445) );
  XNOR2_X1 U560 ( .A(KEYINPUT70), .B(G469), .ZN(n444) );
  XOR2_X1 U561 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n449) );
  NAND2_X1 U562 ( .A1(n446), .A2(G234), .ZN(n447) );
  XNOR2_X1 U563 ( .A(n447), .B(KEYINPUT20), .ZN(n462) );
  NAND2_X1 U564 ( .A1(G217), .A2(n462), .ZN(n448) );
  XNOR2_X1 U565 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U566 ( .A(KEYINPUT25), .B(n450), .ZN(n461) );
  XNOR2_X1 U567 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U568 ( .A(n453), .B(KEYINPUT23), .Z(n455) );
  XNOR2_X1 U569 ( .A(n455), .B(n454), .ZN(n459) );
  NAND2_X1 U570 ( .A1(G234), .A2(n712), .ZN(n457) );
  XOR2_X1 U571 ( .A(KEYINPUT8), .B(n457), .Z(n508) );
  XNOR2_X1 U572 ( .A(n708), .B(n431), .ZN(n458) );
  NOR2_X1 U573 ( .A1(G902), .A2(n691), .ZN(n460) );
  NAND2_X1 U574 ( .A1(n462), .A2(G221), .ZN(n463) );
  XOR2_X1 U575 ( .A(KEYINPUT21), .B(n463), .Z(n648) );
  NAND2_X1 U576 ( .A1(n647), .A2(n648), .ZN(n644) );
  NAND2_X1 U577 ( .A1(n493), .A2(G210), .ZN(n464) );
  XNOR2_X1 U578 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U579 ( .A(n466), .B(KEYINPUT5), .Z(n470) );
  XNOR2_X1 U580 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U582 ( .A(KEYINPUT73), .B(KEYINPUT98), .ZN(n474) );
  NAND2_X1 U583 ( .A1(n476), .A2(G214), .ZN(n477) );
  XNOR2_X1 U584 ( .A(KEYINPUT91), .B(n477), .ZN(n556) );
  INV_X1 U585 ( .A(n556), .ZN(n635) );
  XNOR2_X1 U586 ( .A(n478), .B(KEYINPUT30), .ZN(n488) );
  XNOR2_X1 U587 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U588 ( .A1(G952), .A2(n482), .ZN(n664) );
  NOR2_X1 U589 ( .A1(G953), .A2(n664), .ZN(n564) );
  NOR2_X1 U590 ( .A1(G900), .A2(n562), .ZN(n483) );
  NAND2_X1 U591 ( .A1(G953), .A2(n483), .ZN(n484) );
  XNOR2_X1 U592 ( .A(KEYINPUT107), .B(n484), .ZN(n485) );
  XOR2_X1 U593 ( .A(KEYINPUT82), .B(n486), .Z(n519) );
  XNOR2_X1 U594 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n501) );
  XNOR2_X1 U595 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U596 ( .A(n708), .B(n492), .ZN(n500) );
  NAND2_X1 U597 ( .A1(G214), .A2(n493), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U599 ( .A(n496), .B(G122), .Z(n498) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n500), .B(n499), .ZN(n606) );
  XNOR2_X1 U602 ( .A(n503), .B(n502), .ZN(n507) );
  XNOR2_X1 U603 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U604 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U605 ( .A(n507), .B(n506), .Z(n510) );
  NAND2_X1 U606 ( .A1(G217), .A2(n508), .ZN(n509) );
  XNOR2_X1 U607 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U608 ( .A(n512), .B(n511), .ZN(n602) );
  NOR2_X1 U609 ( .A1(n602), .A2(G902), .ZN(n513) );
  XOR2_X1 U610 ( .A(n513), .B(G478), .Z(n541) );
  INV_X1 U611 ( .A(n541), .ZN(n518) );
  NOR2_X1 U612 ( .A1(n542), .A2(n518), .ZN(n514) );
  XNOR2_X1 U613 ( .A(n514), .B(KEYINPUT106), .ZN(n586) );
  NAND2_X1 U614 ( .A1(n525), .A2(n586), .ZN(n515) );
  NOR2_X1 U615 ( .A1(n516), .A2(n515), .ZN(n621) );
  XOR2_X1 U616 ( .A(KEYINPUT84), .B(n621), .Z(n524) );
  XNOR2_X1 U617 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n517) );
  XOR2_X1 U618 ( .A(KEYINPUT6), .B(n581), .Z(n575) );
  NAND2_X1 U619 ( .A1(n518), .A2(n529), .ZN(n625) );
  INV_X1 U620 ( .A(n625), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n519), .A2(n648), .ZN(n520) );
  NAND2_X1 U622 ( .A1(n527), .A2(n533), .ZN(n521) );
  NAND2_X1 U623 ( .A1(n543), .A2(n554), .ZN(n522) );
  XOR2_X1 U624 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n526) );
  NAND2_X1 U625 ( .A1(n527), .A2(n551), .ZN(n528) );
  XOR2_X1 U626 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n532) );
  XNOR2_X1 U627 ( .A(n530), .B(KEYINPUT104), .ZN(n638) );
  NAND2_X1 U628 ( .A1(n634), .A2(n638), .ZN(n531) );
  XNOR2_X1 U629 ( .A(n532), .B(n531), .ZN(n665) );
  AND2_X1 U630 ( .A1(n651), .A2(n533), .ZN(n534) );
  XNOR2_X1 U631 ( .A(n534), .B(KEYINPUT28), .ZN(n537) );
  NAND2_X1 U632 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U633 ( .A1(n665), .A2(n544), .ZN(n538) );
  XOR2_X1 U634 ( .A(KEYINPUT42), .B(n538), .Z(n722) );
  NAND2_X1 U635 ( .A1(n723), .A2(n722), .ZN(n540) );
  XOR2_X1 U636 ( .A(KEYINPUT46), .B(KEYINPUT86), .Z(n539) );
  XNOR2_X1 U637 ( .A(n540), .B(n539), .ZN(n548) );
  NAND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n628) );
  NAND2_X1 U639 ( .A1(n625), .A2(n628), .ZN(n633) );
  INV_X1 U640 ( .A(n633), .ZN(n545) );
  OR2_X1 U641 ( .A1(n544), .A2(n566), .ZN(n622) );
  NOR2_X1 U642 ( .A1(n545), .A2(n622), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n546), .B(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U644 ( .A1(n548), .A2(n547), .ZN(n549) );
  INV_X1 U645 ( .A(n628), .ZN(n552) );
  NAND2_X1 U646 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n553), .B(KEYINPUT110), .ZN(n724) );
  NAND2_X1 U648 ( .A1(n645), .A2(n554), .ZN(n555) );
  NOR2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U650 ( .A(n557), .B(KEYINPUT43), .ZN(n558) );
  NOR2_X1 U651 ( .A1(n559), .A2(n558), .ZN(n632) );
  XNOR2_X1 U652 ( .A(G898), .B(KEYINPUT93), .ZN(n696) );
  NAND2_X1 U653 ( .A1(n696), .A2(G953), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n561), .B(KEYINPUT94), .ZN(n704) );
  NOR2_X1 U655 ( .A1(n704), .A2(n562), .ZN(n563) );
  NOR2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n614) );
  NOR2_X1 U658 ( .A1(n645), .A2(n644), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n582), .A2(n651), .ZN(n654) );
  XNOR2_X1 U660 ( .A(n569), .B(KEYINPUT31), .ZN(n627) );
  NAND2_X1 U661 ( .A1(n614), .A2(n627), .ZN(n570) );
  AND2_X1 U662 ( .A1(n648), .A2(n638), .ZN(n571) );
  NAND2_X1 U663 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U664 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n573) );
  XNOR2_X1 U665 ( .A(n574), .B(n573), .ZN(n580) );
  INV_X1 U666 ( .A(n575), .ZN(n591) );
  XOR2_X1 U667 ( .A(KEYINPUT79), .B(n591), .Z(n576) );
  NOR2_X1 U668 ( .A1(n647), .A2(n645), .ZN(n577) );
  INV_X1 U669 ( .A(n645), .ZN(n579) );
  NOR2_X1 U670 ( .A1(n580), .A2(n579), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n582), .A2(n591), .ZN(n583) );
  XNOR2_X1 U672 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n647), .A2(n589), .ZN(n590) );
  NOR2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n612) );
  NAND2_X1 U675 ( .A1(n592), .A2(KEYINPUT2), .ZN(n593) );
  XOR2_X1 U676 ( .A(KEYINPUT67), .B(n593), .Z(n594) );
  NAND2_X1 U677 ( .A1(G478), .A2(n347), .ZN(n603) );
  XOR2_X1 U678 ( .A(n606), .B(KEYINPUT59), .Z(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n609) );
  INV_X1 U680 ( .A(KEYINPUT121), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT60), .ZN(n611) );
  XOR2_X1 U682 ( .A(G101), .B(n612), .Z(G3) );
  NOR2_X1 U683 ( .A1(n625), .A2(n614), .ZN(n613) );
  XOR2_X1 U684 ( .A(G104), .B(n613), .Z(G6) );
  NOR2_X1 U685 ( .A1(n628), .A2(n614), .ZN(n616) );
  XNOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(G107), .B(n617), .ZN(G9) );
  XNOR2_X1 U689 ( .A(G110), .B(n618), .ZN(G12) );
  NOR2_X1 U690 ( .A1(n628), .A2(n622), .ZN(n620) );
  XNOR2_X1 U691 ( .A(G128), .B(KEYINPUT29), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(G30) );
  XOR2_X1 U693 ( .A(G143), .B(n621), .Z(G45) );
  NOR2_X1 U694 ( .A1(n625), .A2(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(G146), .B(KEYINPUT111), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(G48) );
  NOR2_X1 U697 ( .A1(n625), .A2(n627), .ZN(n626) );
  XOR2_X1 U698 ( .A(G113), .B(n626), .Z(G15) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U700 ( .A(G116), .B(n629), .Z(G18) );
  XNOR2_X1 U701 ( .A(G125), .B(n630), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n631), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U703 ( .A(G140), .B(n632), .Z(G42) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n641) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT113), .B(n637), .ZN(n639) );
  NAND2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U709 ( .A(KEYINPUT114), .B(n642), .Z(n643) );
  NOR2_X1 U710 ( .A1(n666), .A2(n643), .ZN(n660) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n646), .B(KEYINPUT50), .ZN(n653) );
  NOR2_X1 U713 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(n649), .Z(n650) );
  NOR2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U716 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U717 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U718 ( .A(n656), .B(KEYINPUT112), .ZN(n657) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(n657), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n665), .A2(n658), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U722 ( .A(KEYINPUT115), .B(n661), .Z(n662) );
  XNOR2_X1 U723 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  NOR2_X1 U724 ( .A1(n664), .A2(n663), .ZN(n669) );
  OR2_X1 U725 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U726 ( .A(KEYINPUT116), .B(n667), .Z(n668) );
  NOR2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n670), .A2(n712), .ZN(n678) );
  XNOR2_X1 U729 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n672) );
  NAND2_X1 U730 ( .A1(n697), .A2(n672), .ZN(n671) );
  XNOR2_X1 U731 ( .A(KEYINPUT85), .B(n671), .ZN(n676) );
  NAND2_X1 U732 ( .A1(n672), .A2(n711), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U734 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U736 ( .A(KEYINPUT53), .B(n679), .ZN(G75) );
  XNOR2_X1 U737 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n682) );
  XNOR2_X1 U738 ( .A(n680), .B(KEYINPUT117), .ZN(n681) );
  XNOR2_X1 U739 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT118), .ZN(n684) );
  XOR2_X1 U741 ( .A(n684), .B(KEYINPUT57), .Z(n687) );
  XNOR2_X1 U742 ( .A(n685), .B(KEYINPUT58), .ZN(n686) );
  NOR2_X1 U743 ( .A1(n693), .A2(n689), .ZN(G54) );
  NAND2_X1 U744 ( .A1(G217), .A2(n347), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U746 ( .A1(n693), .A2(n692), .ZN(G66) );
  NAND2_X1 U747 ( .A1(G953), .A2(G224), .ZN(n694) );
  XOR2_X1 U748 ( .A(KEYINPUT61), .B(n694), .Z(n695) );
  NOR2_X1 U749 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U750 ( .A1(G953), .A2(n697), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n699), .A2(n698), .ZN(n706) );
  XNOR2_X1 U752 ( .A(n700), .B(G101), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U755 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U756 ( .A(KEYINPUT124), .B(n707), .ZN(G69) );
  XOR2_X1 U757 ( .A(n709), .B(n708), .Z(n710) );
  XNOR2_X1 U758 ( .A(KEYINPUT125), .B(n710), .ZN(n715) );
  XNOR2_X1 U759 ( .A(n715), .B(n711), .ZN(n713) );
  NAND2_X1 U760 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U761 ( .A(n714), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U762 ( .A(G227), .B(n715), .ZN(n716) );
  NAND2_X1 U763 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U764 ( .A1(G953), .A2(n717), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n719), .A2(n718), .ZN(G72) );
  XNOR2_X1 U766 ( .A(G119), .B(n720), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(KEYINPUT127), .ZN(G21) );
  XNOR2_X1 U768 ( .A(G137), .B(n722), .ZN(G39) );
  XNOR2_X1 U769 ( .A(G131), .B(n723), .ZN(G33) );
  XNOR2_X1 U770 ( .A(G134), .B(n724), .ZN(G36) );
  XNOR2_X1 U771 ( .A(n725), .B(G122), .ZN(G24) );
endmodule

