

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U322 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n511) );
  XNOR2_X1 U324 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U325 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n515) );
  XNOR2_X1 U326 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n516), .B(n515), .ZN(n548) );
  AND2_X1 U328 ( .A1(n557), .A2(n556), .ZN(n568) );
  XOR2_X1 U329 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n291) );
  XNOR2_X1 U330 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n290) );
  XNOR2_X1 U331 ( .A(n291), .B(n290), .ZN(n305) );
  XOR2_X1 U332 ( .A(G155GAT), .B(G162GAT), .Z(n293) );
  XNOR2_X1 U333 ( .A(G120GAT), .B(G148GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U335 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U336 ( .A(G1GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(n297), .B(n296), .Z(n303) );
  XNOR2_X1 U339 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n298), .B(KEYINPUT2), .ZN(n391) );
  XOR2_X1 U341 ( .A(G85GAT), .B(n391), .Z(n300) );
  NAND2_X1 U342 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U344 ( .A(G29GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U346 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U347 ( .A(KEYINPUT83), .B(G134GAT), .Z(n307) );
  XNOR2_X1 U348 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(n308), .ZN(n367) );
  XNOR2_X1 U351 ( .A(n309), .B(n367), .ZN(n552) );
  INV_X1 U352 ( .A(n552), .ZN(n495) );
  XOR2_X1 U353 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n311) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G29GAT), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U356 ( .A(KEYINPUT68), .B(n312), .ZN(n415) );
  XOR2_X1 U357 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n313) );
  XOR2_X1 U359 ( .A(n314), .B(n313), .Z(n328) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G141GAT), .Z(n316) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G113GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U363 ( .A(KEYINPUT70), .B(KEYINPUT65), .Z(n318) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(G8GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U366 ( .A(n320), .B(n319), .Z(n326) );
  XNOR2_X1 U367 ( .A(G15GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n321), .B(KEYINPUT69), .ZN(n436) );
  XOR2_X1 U369 ( .A(G50GAT), .B(n436), .Z(n323) );
  NAND2_X1 U370 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(n324), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n415), .B(n329), .ZN(n574) );
  XNOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n330) );
  XNOR2_X1 U377 ( .A(n330), .B(KEYINPUT71), .ZN(n433) );
  INV_X1 U378 ( .A(n433), .ZN(n331) );
  XOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .Z(n417) );
  NAND2_X1 U380 ( .A1(n331), .A2(n417), .ZN(n334) );
  INV_X1 U381 ( .A(n417), .ZN(n332) );
  NAND2_X1 U382 ( .A1(n433), .A2(n332), .ZN(n333) );
  NAND2_X1 U383 ( .A1(n334), .A2(n333), .ZN(n336) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U386 ( .A(G120GAT), .B(G71GAT), .Z(n351) );
  XNOR2_X1 U387 ( .A(n351), .B(G204GAT), .ZN(n338) );
  INV_X1 U388 ( .A(KEYINPUT73), .ZN(n337) );
  XOR2_X1 U389 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n342) );
  XNOR2_X1 U390 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n341) );
  XOR2_X1 U391 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U392 ( .A(n344), .B(n343), .ZN(n348) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U394 ( .A(n345), .B(G148GAT), .ZN(n393) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n346), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U397 ( .A(n393), .B(n379), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n481) );
  NOR2_X1 U399 ( .A1(n574), .A2(n481), .ZN(n466) );
  XOR2_X1 U400 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n350) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n380) );
  XOR2_X1 U403 ( .A(n351), .B(n380), .Z(n353) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(G99GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n366) );
  XOR2_X1 U406 ( .A(G183GAT), .B(G176GAT), .Z(n355) );
  XNOR2_X1 U407 ( .A(G15GAT), .B(G190GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U409 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n357) );
  XNOR2_X1 U410 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U413 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n361) );
  NAND2_X1 U414 ( .A1(G227GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(KEYINPUT89), .B(n362), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n521) );
  INV_X1 U420 ( .A(n521), .ZN(n556) );
  XOR2_X1 U421 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n373) );
  XOR2_X1 U422 ( .A(G211GAT), .B(G218GAT), .Z(n370) );
  XNOR2_X1 U423 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(G197GAT), .B(n371), .Z(n394) );
  XOR2_X1 U426 ( .A(G8GAT), .B(G183GAT), .Z(n442) );
  XNOR2_X1 U427 ( .A(n394), .B(n442), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n378) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G190GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(KEYINPUT78), .ZN(n425) );
  XOR2_X1 U431 ( .A(n425), .B(KEYINPUT95), .Z(n376) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n378), .B(n377), .Z(n382) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n549) );
  XOR2_X1 U437 ( .A(n549), .B(KEYINPUT27), .Z(n403) );
  NAND2_X1 U438 ( .A1(n403), .A2(n552), .ZN(n517) );
  NOR2_X1 U439 ( .A1(n556), .A2(n517), .ZN(n397) );
  XOR2_X1 U440 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n384) );
  XNOR2_X1 U441 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U443 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n386) );
  XOR2_X1 U444 ( .A(G50GAT), .B(G162GAT), .Z(n416) );
  XOR2_X1 U445 ( .A(G22GAT), .B(G155GAT), .Z(n437) );
  XNOR2_X1 U446 ( .A(n416), .B(n437), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U448 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U451 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n554) );
  XNOR2_X1 U454 ( .A(n554), .B(KEYINPUT28), .ZN(n519) );
  NAND2_X1 U455 ( .A1(n397), .A2(n519), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n398), .B(KEYINPUT98), .ZN(n408) );
  INV_X1 U457 ( .A(n549), .ZN(n472) );
  NAND2_X1 U458 ( .A1(n472), .A2(n556), .ZN(n399) );
  NAND2_X1 U459 ( .A1(n399), .A2(n554), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(KEYINPUT25), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n401), .B(KEYINPUT99), .ZN(n405) );
  NOR2_X1 U462 ( .A1(n554), .A2(n556), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n402), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U464 ( .A1(n403), .A2(n572), .ZN(n404) );
  NAND2_X1 U465 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U466 ( .A1(n495), .A2(n406), .ZN(n407) );
  NAND2_X1 U467 ( .A1(n408), .A2(n407), .ZN(n461) );
  XOR2_X1 U468 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n410) );
  XNOR2_X1 U469 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U471 ( .A(KEYINPUT77), .B(KEYINPUT74), .Z(n412) );
  XNOR2_X1 U472 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n429) );
  INV_X1 U475 ( .A(n415), .ZN(n421) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n419) );
  XNOR2_X1 U477 ( .A(G218GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U480 ( .A1(G232GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(n424), .B(KEYINPUT75), .Z(n427) );
  XNOR2_X1 U483 ( .A(n425), .B(KEYINPUT76), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n546) );
  XOR2_X1 U486 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n435) );
  XOR2_X1 U487 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n431) );
  XNOR2_X1 U488 ( .A(KEYINPUT82), .B(KEYINPUT80), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n449) );
  XOR2_X1 U492 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U493 ( .A1(G231GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n447) );
  XOR2_X1 U495 ( .A(KEYINPUT79), .B(G64GAT), .Z(n441) );
  XNOR2_X1 U496 ( .A(G211GAT), .B(G78GAT), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U498 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U499 ( .A(G127GAT), .B(G71GAT), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n542) );
  INV_X1 U503 ( .A(n542), .ZN(n580) );
  NAND2_X1 U504 ( .A1(n546), .A2(n580), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT16), .B(n450), .Z(n451) );
  AND2_X1 U506 ( .A1(n461), .A2(n451), .ZN(n482) );
  NAND2_X1 U507 ( .A1(n466), .A2(n482), .ZN(n459) );
  NOR2_X1 U508 ( .A1(n495), .A2(n459), .ZN(n453) );
  XNOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U511 ( .A(G1GAT), .B(n454), .Z(G1324GAT) );
  NOR2_X1 U512 ( .A1(n549), .A2(n459), .ZN(n456) );
  XNOR2_X1 U513 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(G1325GAT) );
  NOR2_X1 U515 ( .A1(n521), .A2(n459), .ZN(n458) );
  XNOR2_X1 U516 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(G1326GAT) );
  NOR2_X1 U518 ( .A1(n519), .A2(n459), .ZN(n460) );
  XOR2_X1 U519 ( .A(G22GAT), .B(n460), .Z(G1327GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n468) );
  XNOR2_X1 U521 ( .A(KEYINPUT36), .B(n546), .ZN(n584) );
  NAND2_X1 U522 ( .A1(n542), .A2(n461), .ZN(n462) );
  XNOR2_X1 U523 ( .A(KEYINPUT102), .B(n462), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n584), .A2(n463), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n465), .B(n464), .ZN(n494) );
  NAND2_X1 U527 ( .A1(n466), .A2(n494), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n478) );
  NAND2_X1 U529 ( .A1(n552), .A2(n478), .ZN(n471) );
  XNOR2_X1 U530 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT39), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(G1328GAT) );
  NAND2_X1 U533 ( .A1(n472), .A2(n478), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n475) );
  NAND2_X1 U536 ( .A1(n478), .A2(n556), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U538 ( .A(G43GAT), .B(n476), .Z(G1330GAT) );
  XOR2_X1 U539 ( .A(G50GAT), .B(KEYINPUT107), .Z(n480) );
  INV_X1 U540 ( .A(n519), .ZN(n477) );
  NAND2_X1 U541 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(G1331GAT) );
  INV_X1 U543 ( .A(n574), .ZN(n558) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT41), .ZN(n536) );
  NOR2_X1 U545 ( .A1(n558), .A2(n536), .ZN(n493) );
  NAND2_X1 U546 ( .A1(n493), .A2(n482), .ZN(n489) );
  NOR2_X1 U547 ( .A1(n495), .A2(n489), .ZN(n484) );
  XNOR2_X1 U548 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U550 ( .A(G57GAT), .B(n485), .Z(G1332GAT) );
  NOR2_X1 U551 ( .A1(n549), .A2(n489), .ZN(n487) );
  XNOR2_X1 U552 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(G1333GAT) );
  NOR2_X1 U554 ( .A1(n521), .A2(n489), .ZN(n488) );
  XOR2_X1 U555 ( .A(G71GAT), .B(n488), .Z(G1334GAT) );
  NOR2_X1 U556 ( .A1(n519), .A2(n489), .ZN(n491) );
  XNOR2_X1 U557 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U559 ( .A(G78GAT), .B(n492), .ZN(G1335GAT) );
  NAND2_X1 U560 ( .A1(n494), .A2(n493), .ZN(n501) );
  NOR2_X1 U561 ( .A1(n495), .A2(n501), .ZN(n497) );
  XNOR2_X1 U562 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1336GAT) );
  NOR2_X1 U564 ( .A1(n549), .A2(n501), .ZN(n498) );
  XOR2_X1 U565 ( .A(KEYINPUT112), .B(n498), .Z(n499) );
  XNOR2_X1 U566 ( .A(G92GAT), .B(n499), .ZN(G1337GAT) );
  NOR2_X1 U567 ( .A1(n521), .A2(n501), .ZN(n500) );
  XOR2_X1 U568 ( .A(G99GAT), .B(n500), .Z(G1338GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n501), .ZN(n502) );
  XOR2_X1 U570 ( .A(KEYINPUT44), .B(n502), .Z(n503) );
  XNOR2_X1 U571 ( .A(G106GAT), .B(n503), .ZN(G1339GAT) );
  NOR2_X1 U572 ( .A1(n584), .A2(n542), .ZN(n504) );
  XOR2_X1 U573 ( .A(KEYINPUT45), .B(n504), .Z(n505) );
  NOR2_X1 U574 ( .A1(n481), .A2(n505), .ZN(n506) );
  NAND2_X1 U575 ( .A1(n506), .A2(n574), .ZN(n514) );
  INV_X1 U576 ( .A(n546), .ZN(n569) );
  NOR2_X1 U577 ( .A1(n574), .A2(n536), .ZN(n507) );
  XNOR2_X1 U578 ( .A(n507), .B(KEYINPUT46), .ZN(n508) );
  NOR2_X1 U579 ( .A1(n508), .A2(n580), .ZN(n509) );
  XNOR2_X1 U580 ( .A(n509), .B(KEYINPUT113), .ZN(n510) );
  NOR2_X1 U581 ( .A1(n569), .A2(n510), .ZN(n512) );
  NAND2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n516) );
  NOR2_X1 U583 ( .A1(n517), .A2(n548), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT116), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n533), .A2(n519), .ZN(n520) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n558), .A2(n529), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n524) );
  INV_X1 U590 ( .A(n536), .ZN(n561) );
  NAND2_X1 U591 ( .A1(n529), .A2(n561), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n526) );
  NAND2_X1 U595 ( .A1(n529), .A2(n580), .ZN(n525) );
  XNOR2_X1 U596 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n531) );
  NAND2_X1 U599 ( .A1(n529), .A2(n569), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  NAND2_X1 U602 ( .A1(n572), .A2(n533), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n574), .A2(n545), .ZN(n534) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n534), .Z(n535) );
  XNOR2_X1 U605 ( .A(KEYINPUT120), .B(n535), .ZN(G1344GAT) );
  NOR2_X1 U606 ( .A1(n536), .A2(n545), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n538) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n537) );
  XNOR2_X1 U609 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(KEYINPUT53), .B(n539), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n542), .A2(n545), .ZN(n544) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(KEYINPUT123), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n547), .Z(G1347GAT) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U619 ( .A(KEYINPUT54), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n573) );
  NAND2_X1 U622 ( .A1(n573), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(KEYINPUT55), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n568), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT125), .Z(n563) );
  NAND2_X1 U627 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n568), .A2(n580), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT126), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(n567), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n571), .ZN(G1351GAT) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n583) );
  NOR2_X1 U638 ( .A1(n574), .A2(n583), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U643 ( .A(n583), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n581), .A2(n481), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

