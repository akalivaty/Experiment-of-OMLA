//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT74), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(KEYINPUT23), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT64), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(G169gat), .C2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT65), .B(G183gat), .Z(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT24), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n219), .A2(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT25), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n222), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n220), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT25), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n217), .A3(new_n212), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT27), .ZN(new_n234));
  AOI21_X1  g033(.A(G190gat), .B1(new_n234), .B2(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT28), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT66), .B1(new_n219), .B2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n219), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n235), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n223), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n245), .B1(KEYINPUT26), .B2(new_n211), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n210), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n233), .B(KEYINPUT72), .C1(new_n244), .C2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n235), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n243), .B1(new_n251), .B2(new_n239), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(new_n237), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n253), .B2(new_n232), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  AOI211_X1 g057(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT69), .B(G120gat), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n260), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT67), .B(G127gat), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G134gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT1), .B1(new_n257), .B2(new_n258), .ZN(new_n267));
  NAND2_X1  g066(.A1(G113gat), .A2(G120gat), .ZN(new_n268));
  INV_X1    g067(.A(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(G134gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n266), .B1(new_n265), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n272), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT71), .A3(new_n263), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n249), .A2(new_n254), .A3(new_n277), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n280), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n253), .A2(new_n232), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT72), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n207), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(KEYINPUT73), .B1(KEYINPUT32), .B2(new_n287), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n207), .A2(new_n288), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n281), .A2(new_n286), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(new_n282), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n283), .B1(new_n281), .B2(new_n286), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT75), .A2(KEYINPUT34), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n290), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n298), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(KEYINPUT73), .A3(new_n206), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n293), .A3(new_n206), .ZN(new_n308));
  INV_X1    g107(.A(new_n292), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n303), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n202), .B1(new_n301), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n300), .B1(new_n290), .B2(new_n294), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n310), .A3(new_n303), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT36), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  AND2_X1   g116(.A1(G211gat), .A2(G218gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(KEYINPUT22), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G211gat), .B(G218gat), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G148gat), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(G141gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT79), .B(G141gat), .Z(new_n335));
  OAI21_X1  g134(.A(new_n324), .B1(new_n335), .B2(new_n322), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n327), .B1(new_n332), .B2(KEYINPUT2), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n321), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n321), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n344));
  INV_X1    g143(.A(new_n338), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G78gat), .B(G106gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G22gat), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT31), .B(G50gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n348), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n275), .A3(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n277), .A2(new_n280), .A3(new_n338), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n345), .B2(new_n275), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n279), .A2(KEYINPUT81), .A3(new_n338), .A4(new_n263), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n355), .B(new_n358), .C1(new_n361), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n355), .A2(new_n356), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(new_n360), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n362), .A3(new_n365), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n364), .A2(new_n365), .B1(new_n345), .B2(new_n275), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT5), .B1(new_n372), .B2(new_n356), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT0), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n367), .B(new_n378), .C1(new_n371), .C2(new_n373), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT82), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n380), .A2(new_n385), .A3(new_n381), .A4(new_n382), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n379), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G226gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT29), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n233), .B(new_n394), .C1(new_n244), .C2(new_n248), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT76), .B1(new_n253), .B2(new_n232), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n285), .A2(new_n391), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n321), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n391), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n253), .B2(new_n232), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n343), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n402), .A4(new_n406), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT77), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n402), .A3(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT77), .B1(new_n408), .B2(new_n409), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n353), .B1(new_n388), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n316), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n355), .B1(new_n361), .B2(new_n366), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n357), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT39), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n372), .B2(new_n356), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n421), .A3(new_n357), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n424), .A2(KEYINPUT83), .A3(new_n378), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT83), .B1(new_n424), .B2(new_n378), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT40), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n408), .A3(new_n409), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n429), .A2(new_n380), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n383), .A2(new_n387), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n407), .B1(new_n403), .B2(KEYINPUT37), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n399), .B2(new_n402), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT38), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT84), .B(KEYINPUT38), .C1(new_n434), .C2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(new_n411), .ZN(new_n441));
  INV_X1    g240(.A(new_n434), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n400), .A2(new_n321), .A3(new_n401), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n443), .A2(KEYINPUT37), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n343), .B1(new_n397), .B2(new_n398), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT38), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n433), .A2(new_n439), .A3(new_n440), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n448), .A3(new_n353), .ZN(new_n449));
  INV_X1    g248(.A(new_n353), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n313), .B2(new_n314), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n388), .A3(new_n416), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT85), .B1(new_n433), .B2(new_n431), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n383), .A2(new_n387), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456));
  INV_X1    g255(.A(new_n431), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n451), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n418), .A2(new_n449), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n462));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G1gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT16), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n463), .ZN(new_n468));
  INV_X1    g267(.A(G8gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n464), .A3(G1gat), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT15), .ZN(new_n474));
  NOR2_X1   g273(.A1(G43gat), .A2(G50gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G43gat), .A2(G50gat), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(new_n475), .A3(KEYINPUT15), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G29gat), .A2(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT88), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n482), .A2(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT15), .B1(new_n479), .B2(new_n475), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n482), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n490), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n478), .ZN(new_n498));
  AOI221_X4 g297(.A(KEYINPUT17), .B1(new_n481), .B2(new_n491), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n498), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n491), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n462), .B(new_n473), .C1(new_n499), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n466), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n463), .A2(new_n467), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n470), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G8gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n502), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT17), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n494), .A2(new_n498), .B1(new_n491), .B2(new_n481), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n500), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT91), .B1(new_n473), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n504), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT18), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n518), .B(KEYINPUT13), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n473), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n510), .A2(new_n511), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT11), .B(G169gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT18), .B1(new_n517), .B2(new_n518), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n526), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n518), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n473), .B1(new_n499), .B2(new_n503), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n462), .B1(new_n510), .B2(new_n511), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n539), .B2(new_n504), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n524), .B1(new_n540), .B2(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n518), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n532), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n535), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n461), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G190gat), .B(G218gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT101), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT41), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT98), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  INV_X1    g359(.A(new_n558), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(G92gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(KEYINPUT8), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n563), .A2(new_n569), .A3(new_n567), .A4(new_n570), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n564), .A2(new_n571), .A3(KEYINPUT99), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n555), .B1(new_n577), .B2(new_n511), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT100), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n576), .B(new_n575), .C1(new_n499), .C2(new_n503), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n554), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n552), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n582), .A3(new_n551), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n330), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT93), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n595), .A2(new_n596), .A3(new_n600), .A4(new_n597), .ZN(new_n601));
  NOR2_X1   g400(.A1(G57gat), .A2(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604));
  NAND2_X1  g403(.A1(G57gat), .A2(G64gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT94), .B1(new_n607), .B2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n599), .B(new_n601), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n593), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n603), .A3(new_n605), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n613), .A2(KEYINPUT96), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT96), .B1(new_n613), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n510), .B1(new_n619), .B2(KEYINPUT21), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n613), .A2(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n624), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G127gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n624), .B(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n269), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n621), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n630), .A3(new_n621), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n592), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n592), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n588), .A2(new_n637), .A3(KEYINPUT102), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n585), .A2(new_n587), .ZN(new_n640));
  INV_X1    g439(.A(new_n633), .ZN(new_n641));
  INV_X1    g440(.A(new_n592), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n641), .A2(new_n631), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n639), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n613), .A2(new_n572), .A3(new_n616), .A4(new_n574), .ZN(new_n648));
  INV_X1    g447(.A(new_n622), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n647), .B(new_n648), .C1(new_n577), .C2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n613), .A2(KEYINPUT96), .A3(new_n616), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n577), .A2(new_n652), .A3(KEYINPUT10), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT103), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n648), .B1(new_n577), .B2(new_n649), .ZN(new_n660));
  INV_X1    g459(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n666), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n661), .B1(new_n650), .B2(new_n654), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n547), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n388), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n466), .ZN(G1324gat));
  AND2_X1   g477(.A1(new_n312), .A2(new_n315), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n388), .A2(new_n416), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n450), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n449), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n453), .A2(new_n460), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n546), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n431), .A3(new_n685), .A4(new_n675), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G8gat), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT16), .B(G8gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT105), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n688), .B2(new_n689), .ZN(new_n695));
  OAI221_X1 g494(.A(new_n690), .B1(new_n686), .B2(new_n694), .C1(new_n695), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g495(.A(G15gat), .B1(new_n676), .B2(new_n679), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n301), .A2(new_n311), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n676), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n676), .A2(new_n353), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n388), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n644), .A2(new_n674), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n588), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n547), .A2(new_n484), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n461), .B2(new_n588), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n640), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT106), .B1(new_n535), .B2(new_n545), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n535), .A2(new_n545), .A3(KEYINPUT106), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n705), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n712), .A2(new_n704), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n708), .B1(new_n484), .B2(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  AOI211_X1 g520(.A(G36gat), .B(new_n457), .C1(new_n721), .C2(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n547), .A2(new_n706), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n712), .A2(new_n431), .A3(new_n718), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n485), .ZN(G1329gat));
  NOR2_X1   g526(.A1(new_n698), .A2(G43gat), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n684), .A2(new_n685), .A3(new_n706), .A4(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n711), .A3(new_n316), .A4(new_n718), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(G43gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g531(.A1(new_n684), .A2(new_n450), .A3(new_n685), .A4(new_n706), .ZN(new_n733));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(KEYINPUT48), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n353), .A2(new_n734), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n710), .A2(new_n711), .A3(new_n718), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1331gat));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n638), .B(new_n645), .C1(new_n714), .C2(new_n715), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n674), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n461), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n684), .A2(KEYINPUT109), .A3(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n704), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g550(.A(KEYINPUT49), .B(G64gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n431), .A3(new_n752), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n748), .A2(new_n457), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n748), .B2(new_n679), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n698), .A2(G71gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n746), .A2(new_n747), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(KEYINPUT50), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n749), .A2(new_n450), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g564(.A(new_n588), .B1(new_n682), .B2(new_n683), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n716), .A2(new_n637), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(new_n566), .A3(new_n704), .A4(new_n673), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n716), .A2(new_n637), .A3(new_n674), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n712), .A2(new_n704), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n775), .B2(new_n566), .ZN(G1336gat));
  NAND4_X1  g575(.A1(new_n710), .A2(new_n711), .A3(new_n431), .A4(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(new_n565), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n457), .A2(G92gat), .A3(new_n674), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n771), .B1(new_n766), .B2(new_n767), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n780), .B(KEYINPUT111), .Z(new_n786));
  AOI22_X1  g585(.A1(new_n772), .A2(new_n786), .B1(new_n777), .B2(new_n778), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n784), .ZN(G1337gat));
  NOR2_X1   g587(.A1(new_n698), .A2(G99gat), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n673), .B(new_n789), .C1(new_n781), .C2(new_n782), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n710), .A2(new_n711), .A3(new_n316), .A4(new_n774), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G99gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  NOR2_X1   g596(.A1(new_n353), .A2(G106gat), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n673), .B(new_n798), .C1(new_n781), .C2(new_n782), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n710), .A2(new_n711), .A3(new_n450), .A4(new_n774), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n667), .B1(new_n659), .B2(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n650), .A2(new_n654), .A3(new_n657), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT54), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n670), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n647), .B1(new_n575), .B2(new_n576), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n658), .B1(new_n619), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n650), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n655), .A2(new_n656), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n807), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n657), .B1(new_n650), .B2(new_n654), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n666), .B1(new_n819), .B2(new_n813), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n671), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n812), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT55), .B1(new_n810), .B2(new_n670), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n822), .B(new_n672), .C1(new_n824), .C2(new_n808), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n715), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n672), .B1(new_n824), .B2(new_n808), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n825), .A4(new_n812), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n827), .A2(new_n828), .A3(new_n713), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n541), .A2(new_n532), .A3(new_n544), .ZN(new_n834));
  INV_X1    g633(.A(new_n530), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n522), .A2(new_n523), .A3(new_n521), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT115), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n539), .A2(new_n536), .A3(new_n504), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n673), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n640), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n640), .A2(new_n834), .A3(new_n840), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n827), .A3(new_n832), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n644), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n743), .A2(new_n673), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n451), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n388), .A2(new_n431), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n546), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n853), .B(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n716), .A2(new_n257), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n673), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(G120gat), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT117), .B(new_n258), .C1(new_n853), .C2(new_n673), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n673), .A2(new_n262), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n861), .A2(new_n862), .B1(new_n856), .B2(new_n863), .ZN(G1341gat));
  NAND2_X1  g663(.A1(new_n853), .A2(new_n637), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n264), .ZN(G1342gat));
  AND2_X1   g665(.A1(new_n849), .A2(new_n451), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(new_n270), .A3(new_n640), .A4(new_n851), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n868), .B2(KEYINPUT56), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n588), .A3(new_n852), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n270), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n870), .A2(new_n270), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n679), .A2(new_n851), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n679), .A2(KEYINPUT119), .A3(new_n851), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n353), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n808), .B2(new_n811), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n821), .B(new_n886), .C1(new_n535), .C2(new_n545), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(KEYINPUT121), .A3(new_n841), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT121), .B1(new_n887), .B2(new_n841), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n588), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n637), .B1(new_n890), .B2(new_n844), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(new_n847), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT122), .B(new_n884), .C1(new_n891), .C2(new_n847), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(new_n849), .B2(new_n450), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n685), .B(new_n882), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n335), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n849), .A2(new_n450), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n900), .A2(G141gat), .A3(new_n546), .A4(new_n878), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n716), .B(new_n882), .C1(new_n896), .C2(new_n897), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n335), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n322), .A2(KEYINPUT59), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n882), .B1(new_n896), .B2(new_n897), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n674), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n674), .B1(new_n880), .B2(new_n881), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n646), .A2(new_n546), .A3(new_n674), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n843), .A2(new_n825), .A3(new_n812), .A4(new_n830), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n637), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n883), .B(new_n450), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n353), .B1(new_n846), .B2(new_n848), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n911), .B(new_n915), .C1(new_n916), .C2(new_n883), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT59), .B1(new_n918), .B2(new_n322), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n900), .A2(new_n878), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n322), .A3(new_n673), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n909), .B2(new_n644), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n330), .A3(new_n637), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n909), .B2(new_n588), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n331), .A3(new_n640), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n704), .A2(new_n457), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n849), .A2(new_n451), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n716), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n546), .A2(new_n208), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(G1348gat));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n673), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(G176gat), .ZN(G1349gat));
  XNOR2_X1  g735(.A(KEYINPUT27), .B(G183gat), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n931), .A2(new_n637), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n219), .B1(new_n931), .B2(new_n637), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT60), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT60), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1350gat));
  NAND4_X1  g741(.A1(new_n849), .A2(new_n451), .A3(new_n640), .A4(new_n930), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(G190gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(G190gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1351gat));
  XNOR2_X1  g751(.A(KEYINPUT124), .B(G197gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n316), .A2(new_n704), .A3(new_n457), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n915), .B(new_n954), .C1(new_n916), .C2(new_n883), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(new_n546), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n916), .A2(new_n954), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n717), .A2(new_n953), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(new_n957), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n674), .A2(G204gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  OAI21_X1  g762(.A(G204gat), .B1(new_n955), .B2(new_n674), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n962), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT125), .B1(new_n962), .B2(KEYINPUT62), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n963), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n960), .A2(new_n968), .A3(new_n637), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n972), .A2(new_n637), .A3(new_n915), .A4(new_n954), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(KEYINPUT126), .B2(new_n970), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n974), .B(new_n971), .C1(new_n955), .C2(new_n644), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n969), .B1(new_n975), .B2(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n955), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n640), .B1(new_n955), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g780(.A(G218gat), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n588), .A2(G218gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n982), .B1(new_n957), .B2(new_n983), .ZN(G1355gat));
endmodule


