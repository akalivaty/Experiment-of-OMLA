//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT64), .Z(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n210), .B(new_n214), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G68), .B(G77), .ZN(new_n233));
  INV_X1    g0033(.A(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT66), .B(G50), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(KEYINPUT84), .ZN(new_n242));
  INV_X1    g0042(.A(G1), .ZN(new_n243));
  OAI21_X1  g0043(.A(new_n243), .B1(G41), .B2(G45), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n207), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G232), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n249), .A2(new_n248), .ZN(new_n255));
  INV_X1    g0055(.A(new_n207), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(new_n251), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT81), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G87), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1698), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n264), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G226), .A2(G1698), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT80), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT76), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G33), .ZN(new_n278));
  AND4_X1   g0078(.A1(KEYINPUT80), .A2(new_n278), .A3(new_n265), .A4(new_n272), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n261), .B(new_n271), .C1(new_n273), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n256), .A2(new_n249), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n268), .A2(KEYINPUT80), .A3(new_n272), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n265), .A3(new_n272), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT80), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n261), .B1(new_n288), .B2(new_n271), .ZN(new_n289));
  OAI211_X1 g0089(.A(G179), .B(new_n260), .C1(new_n283), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n278), .A2(new_n265), .A3(new_n270), .ZN(new_n291));
  INV_X1    g0091(.A(new_n264), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n284), .B2(new_n287), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n281), .B1(new_n294), .B2(new_n261), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n271), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT81), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n259), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n290), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G58), .A2(G68), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(G20), .B1(new_n302), .B2(new_n201), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G159), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT77), .B(G20), .C1(new_n302), .C2(new_n201), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(G20), .B1(new_n278), .B2(new_n265), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n268), .A2(KEYINPUT7), .A3(G20), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT16), .B(new_n309), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n311), .A2(G20), .ZN(new_n317));
  AOI21_X1  g0117(.A(G33), .B1(new_n275), .B2(new_n277), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n274), .A2(G33), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n311), .B1(new_n322), .B2(G20), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT69), .B1(new_n211), .B2(new_n262), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n328), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n207), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n314), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n243), .A2(G13), .A3(G20), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n243), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n334), .A2(new_n336), .B1(new_n333), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT79), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT79), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n340), .A3(new_n337), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n300), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT18), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n331), .A2(new_n340), .A3(new_n337), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n331), .B2(new_n337), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n300), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n260), .B1(new_n283), .B2(new_n289), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G200), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n331), .A2(new_n337), .ZN(new_n352));
  OAI211_X1 g0152(.A(G190), .B(new_n260), .C1(new_n283), .C2(new_n289), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT82), .A4(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT83), .A4(new_n353), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT82), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n349), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G1698), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n322), .A2(G222), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n322), .A2(G1698), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n364), .B1(new_n365), .B2(new_n322), .C1(new_n366), .C2(new_n269), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n282), .ZN(new_n368));
  INV_X1    g0168(.A(new_n258), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G226), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n253), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(G179), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n306), .A2(G150), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n208), .A2(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n374), .C1(new_n335), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G50), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n330), .B1(new_n377), .B2(new_n333), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n243), .A2(G20), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n334), .A2(G50), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n371), .A2(new_n299), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n372), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT10), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(G200), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(KEYINPUT9), .A3(new_n380), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n368), .A2(G190), .A3(new_n253), .A4(new_n370), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT9), .B1(new_n378), .B2(new_n380), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT73), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n385), .A3(new_n391), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n384), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n306), .A2(G50), .ZN(new_n396));
  XOR2_X1   g0196(.A(new_n396), .B(KEYINPUT74), .Z(new_n397));
  OAI22_X1  g0197(.A1(new_n375), .A2(new_n365), .B1(new_n208), .B2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n330), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT11), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT11), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n330), .C1(new_n397), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n332), .B(KEYINPUT71), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT12), .B1(new_n404), .B2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(G13), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G1), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT12), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G20), .A4(new_n316), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n332), .B(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n330), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n316), .B1(new_n243), .B2(G20), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n405), .A2(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n322), .A2(G226), .A3(new_n363), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n366), .C2(new_n254), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n418), .A2(new_n282), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n257), .A2(G238), .A3(new_n244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n253), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT13), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n253), .A2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n282), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT14), .B1(new_n427), .B2(new_n299), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n426), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n422), .A2(G179), .A3(new_n426), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT75), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n415), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n415), .ZN(new_n436));
  INV_X1    g0236(.A(G190), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n427), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n322), .A2(G232), .A3(new_n363), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  INV_X1    g0244(.A(G238), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n443), .B1(new_n444), .B2(new_n322), .C1(new_n366), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n282), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n369), .A2(G244), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n253), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(G179), .ZN(new_n450));
  INV_X1    g0250(.A(new_n335), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n306), .B1(G20), .B2(G77), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT70), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n375), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n330), .B1(new_n365), .B2(new_n411), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n412), .A2(G77), .A3(new_n379), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT72), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT72), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n412), .A2(new_n460), .A3(G77), .A4(new_n379), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n449), .A2(new_n299), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n450), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n449), .A2(G200), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n447), .A2(G190), .A3(new_n253), .A4(new_n448), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n457), .A3(new_n462), .A4(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n395), .A2(new_n435), .A3(new_n442), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n242), .B1(new_n362), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n435), .A2(new_n442), .ZN(new_n472));
  INV_X1    g0272(.A(new_n394), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n469), .B(new_n383), .C1(new_n473), .C2(new_n392), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n358), .B2(new_n355), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT84), .A4(new_n349), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n333), .A2(new_n444), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT25), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n262), .A2(G1), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n330), .A2(new_n333), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(G107), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT90), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n263), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n278), .A2(new_n208), .A3(new_n265), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n265), .A2(new_n319), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n208), .A2(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n444), .A3(G20), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n493), .A2(KEYINPUT89), .B1(KEYINPUT23), .B2(G107), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n492), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n495), .A2(new_n496), .B1(new_n498), .B2(new_n208), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n488), .A2(new_n491), .A3(new_n494), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT24), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n495), .A2(new_n496), .B1(new_n492), .B2(new_n444), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n493), .A2(KEYINPUT89), .B1(new_n503), .B2(G20), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n488), .A4(new_n491), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n485), .B1(new_n508), .B2(new_n330), .ZN(new_n509));
  INV_X1    g0309(.A(new_n330), .ZN(new_n510));
  AOI211_X1 g0310(.A(KEYINPUT90), .B(new_n510), .C1(new_n501), .C2(new_n507), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n484), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n278), .A2(new_n265), .ZN(new_n513));
  INV_X1    g0313(.A(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G250), .B2(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n513), .A2(new_n516), .B1(new_n262), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n243), .A2(G45), .ZN(new_n519));
  OR2_X1    g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n251), .B2(new_n250), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n518), .A2(new_n282), .B1(new_n523), .B2(G264), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT91), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n257), .A3(G274), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT86), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n252), .A2(new_n528), .A3(new_n522), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n524), .A2(new_n525), .A3(G179), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n518), .A2(new_n282), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n523), .A2(G264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT91), .B1(new_n534), .B2(G169), .ZN(new_n535));
  INV_X1    g0335(.A(G179), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n512), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n444), .B1(new_n321), .B2(new_n323), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n306), .A2(G77), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  INV_X1    g0342(.A(G97), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(G97), .B(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n541), .B1(new_n546), .B2(new_n208), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n330), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n332), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n483), .B2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n527), .A2(new_n529), .B1(new_n523), .B2(G257), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT4), .B1(new_n268), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n322), .A2(G250), .A3(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n553), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(new_n363), .A3(new_n265), .A4(new_n319), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G283), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n282), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n551), .B1(new_n565), .B2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n552), .A2(new_n564), .A3(G190), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n523), .A2(G257), .ZN(new_n568));
  AND4_X1   g0368(.A1(new_n528), .A2(new_n522), .A3(new_n257), .A4(G274), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n528), .B1(new_n252), .B2(new_n522), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n556), .A2(new_n559), .A3(new_n562), .ZN(new_n572));
  INV_X1    g0372(.A(new_n554), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n557), .B1(new_n513), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n281), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G169), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n552), .A2(new_n564), .A3(G179), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n566), .A2(new_n567), .B1(new_n578), .B2(new_n551), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n534), .A2(new_n439), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n534), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n484), .C1(new_n511), .C2(new_n509), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n539), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  INV_X1    g0384(.A(G45), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(G1), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n586), .A2(G250), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n247), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n257), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G238), .A2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n553), .B2(G1698), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n268), .A2(new_n591), .B1(G33), .B2(G116), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n584), .B(new_n589), .C1(new_n592), .C2(new_n281), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n278), .A3(new_n265), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n281), .B1(new_n594), .B2(new_n497), .ZN(new_n595));
  INV_X1    g0395(.A(new_n589), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT87), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n439), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n268), .A2(new_n208), .A3(G68), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n208), .B1(new_n417), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n263), .A2(new_n543), .A3(new_n444), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n330), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n455), .A2(new_n411), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n483), .A2(G87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n593), .A2(new_n597), .A3(G190), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT88), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n593), .A2(new_n597), .A3(new_n612), .A4(G190), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n598), .B(new_n609), .C1(new_n611), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n514), .A2(new_n363), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(G264), .B2(new_n363), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n513), .A2(new_n616), .B1(new_n617), .B2(new_n322), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n282), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n523), .A2(G270), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n530), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(G20), .B1(new_n262), .B2(G97), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n560), .A2(new_n561), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT85), .B1(G33), .B2(G283), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G20), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n330), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT20), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n482), .A2(new_n626), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n510), .A2(new_n404), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n411), .A2(new_n626), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT20), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n330), .A2(new_n625), .A3(new_n633), .A4(new_n627), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n631), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n621), .A2(G169), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n621), .A2(G200), .ZN(new_n639));
  INV_X1    g0439(.A(new_n635), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n618), .A2(new_n282), .B1(new_n523), .B2(G270), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(G190), .A3(new_n530), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n635), .A2(G179), .A3(new_n641), .A4(new_n530), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n621), .A2(KEYINPUT21), .A3(G169), .A4(new_n635), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n638), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n593), .A2(new_n597), .A3(new_n536), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n483), .A2(new_n454), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n606), .A2(new_n648), .A3(new_n607), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n593), .A2(new_n597), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n299), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n614), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n479), .A2(new_n583), .A3(new_n653), .ZN(G372));
  AND3_X1   g0454(.A1(new_n300), .A2(new_n347), .A3(new_n338), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n347), .B1(new_n300), .B2(new_n338), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT75), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n433), .B(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n430), .B1(new_n429), .B2(G169), .ZN(new_n660));
  AOI211_X1 g0460(.A(KEYINPUT14), .B(new_n299), .C1(new_n422), .C2(new_n426), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n436), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n465), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n442), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n356), .A2(new_n357), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n361), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n657), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n393), .A2(new_n394), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n384), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n479), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n645), .A2(new_n644), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n299), .B1(new_n641), .B2(new_n530), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT21), .B1(new_n674), .B2(new_n635), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n539), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n299), .B1(new_n595), .B2(new_n596), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n647), .A2(new_n649), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n611), .A2(new_n613), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n595), .A2(new_n596), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n439), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n609), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n677), .A2(new_n582), .A3(new_n579), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT92), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n576), .A2(new_n688), .A3(new_n577), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n687), .A2(new_n551), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT26), .B1(new_n690), .B2(new_n684), .ZN(new_n691));
  INV_X1    g0491(.A(new_n650), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n593), .A2(new_n597), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(G169), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n598), .A2(new_n609), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n680), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n551), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n576), .B2(new_n577), .ZN(new_n698));
  AND4_X1   g0498(.A1(KEYINPUT26), .A2(new_n694), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n685), .B(new_n686), .C1(new_n691), .C2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n671), .B1(new_n672), .B2(new_n701), .ZN(G369));
  NAND3_X1  g0502(.A1(new_n638), .A2(new_n644), .A3(new_n645), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n407), .A2(new_n208), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(G213), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n640), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n646), .B2(new_n711), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n512), .A2(new_n709), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n539), .A2(new_n717), .A3(new_n582), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n512), .A2(new_n538), .A3(new_n709), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n512), .A2(new_n538), .A3(new_n710), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n703), .A2(new_n710), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n539), .A3(new_n582), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n212), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n602), .A2(G116), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n205), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n552), .A2(new_n524), .A3(new_n564), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n641), .A2(G179), .A3(new_n530), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n693), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT93), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n651), .A2(new_n536), .A3(new_n621), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT30), .A4(new_n734), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n565), .A3(new_n534), .A4(new_n621), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n738), .A2(new_n739), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT31), .B1(new_n745), .B2(new_n709), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n583), .A2(new_n653), .A3(new_n710), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n679), .B(KEYINPUT95), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n680), .A2(new_n683), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n686), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n687), .A2(new_n551), .A3(new_n689), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT26), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT26), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n694), .A2(new_n696), .A3(new_n759), .A4(new_n698), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n685), .A2(new_n754), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n710), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT29), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n700), .A2(new_n764), .A3(new_n710), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n753), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n733), .B1(new_n767), .B2(G1), .ZN(G364));
  NOR2_X1   g0568(.A1(new_n406), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n243), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n728), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n716), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n713), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n207), .B1(G20), .B2(new_n299), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n208), .A2(new_n437), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n536), .A2(G200), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(new_n536), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT33), .B(G317), .Z(new_n789));
  OAI22_X1  g0589(.A1(new_n783), .A2(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n208), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n778), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n489), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n439), .A2(G179), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n777), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(G303), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G179), .A2(G200), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n208), .B1(new_n802), .B2(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n801), .A2(G326), .B1(new_n804), .B2(G294), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n792), .A2(KEYINPUT99), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n792), .A2(KEYINPUT99), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n802), .A3(new_n807), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G283), .A2(new_n809), .B1(new_n811), .B2(G329), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n791), .A2(new_n799), .A3(new_n805), .A4(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n322), .B1(new_n793), .B2(new_n365), .C1(new_n263), .C2(new_n797), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n803), .A2(new_n543), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G50), .B2(new_n801), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n316), .B2(new_n788), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(G107), .C2(new_n809), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT32), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n782), .B(KEYINPUT98), .Z(new_n822));
  OAI211_X1 g0622(.A(new_n818), .B(new_n821), .C1(new_n234), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n776), .B1(new_n813), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G13), .A2(G33), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n775), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n268), .A2(new_n727), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n585), .B2(new_n206), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(KEYINPUT96), .B1(new_n237), .B2(G45), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(KEYINPUT96), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n727), .A2(new_n489), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G355), .B1(new_n626), .B2(new_n727), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n829), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n772), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n824), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n827), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n713), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n774), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  OAI221_X1 g0644(.A(new_n268), .B1(new_n377), .B2(new_n797), .C1(new_n234), .C2(new_n803), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n316), .A2(new_n808), .B1(new_n810), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n793), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n801), .A2(G137), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n788), .C1(new_n822), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n845), .B(new_n847), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n800), .A2(new_n617), .B1(new_n793), .B2(new_n626), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G283), .B2(new_n787), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n809), .A2(G87), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n322), .B(new_n815), .C1(G107), .C2(new_n798), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n782), .A2(G294), .B1(G311), .B2(new_n811), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n776), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n775), .A2(new_n825), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n772), .B1(new_n865), .B2(G77), .ZN(new_n866));
  OR3_X1    g0666(.A1(new_n863), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT102), .B1(new_n863), .B2(new_n866), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n664), .A2(new_n710), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n463), .A2(new_n709), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n468), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n465), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n867), .B(new_n868), .C1(new_n826), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n701), .B2(new_n709), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n469), .A2(new_n710), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n700), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n752), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n839), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n752), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(G384));
  INV_X1    g0684(.A(new_n546), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n209), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT36), .Z(new_n889));
  NOR3_X1   g0689(.A1(new_n205), .A2(new_n365), .A3(new_n302), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n890), .A2(KEYINPUT103), .B1(new_n377), .B2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n243), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n415), .A2(new_n709), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n663), .B2(new_n441), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n435), .A2(new_n442), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n873), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n745), .A2(new_n709), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT31), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n750), .A3(new_n749), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n314), .A2(new_n330), .ZN(new_n905));
  INV_X1    g0705(.A(new_n315), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT7), .B1(new_n268), .B2(G20), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n310), .A2(new_n311), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(G68), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n906), .B1(new_n909), .B2(new_n309), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n337), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n707), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n343), .A2(new_n348), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n668), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n353), .A2(new_n331), .A3(new_n337), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n295), .A2(new_n297), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n439), .B1(new_n918), .B2(new_n260), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n350), .A2(G169), .ZN(new_n921));
  INV_X1    g0721(.A(new_n910), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n330), .A3(new_n314), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n921), .A2(new_n290), .B1(new_n923), .B2(new_n337), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n342), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n346), .A2(KEYINPUT106), .A3(new_n300), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n339), .A2(new_n341), .A3(new_n912), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n338), .B1(G190), .B2(new_n298), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT37), .B1(new_n932), .B2(new_n351), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(KEYINPUT105), .B(KEYINPUT37), .C1(new_n920), .C2(new_n924), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n916), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n904), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n300), .A2(new_n338), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n931), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT37), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT107), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n948), .A3(KEYINPUT37), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n934), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n931), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n655), .A2(new_n656), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n668), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n942), .B1(new_n937), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n479), .A2(new_n903), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n959), .A2(new_n715), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n937), .B2(new_n954), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT38), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n913), .B1(new_n477), .B2(new_n349), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n927), .A2(new_n934), .A3(new_n935), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n936), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(KEYINPUT39), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n435), .A2(new_n709), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n657), .A2(new_n912), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n967), .A2(new_n968), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT104), .ZN(new_n975));
  INV_X1    g0775(.A(new_n869), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n700), .B2(new_n878), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n897), .A2(new_n898), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n975), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n700), .A2(new_n878), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n978), .B(KEYINPUT104), .C1(new_n981), .C2(new_n976), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n974), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n971), .A2(new_n973), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n479), .A2(new_n766), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n671), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n984), .B(new_n986), .Z(new_n987));
  OAI22_X1  g0787(.A1(new_n961), .A2(new_n987), .B1(new_n243), .B2(new_n769), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n961), .A2(new_n987), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n894), .B1(new_n988), .B2(new_n989), .ZN(G367));
  NAND2_X1  g0790(.A1(new_n690), .A2(new_n709), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n579), .B1(new_n697), .B2(new_n710), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n725), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT42), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n539), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n710), .B1(new_n996), .B2(new_n698), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n609), .A2(new_n709), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n684), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n679), .A2(new_n609), .A3(new_n709), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n721), .A2(new_n993), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n728), .B(KEYINPUT41), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n991), .A2(new_n992), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(new_n725), .A3(new_n722), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1011), .B1(new_n722), .B2(new_n725), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n721), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(KEYINPUT109), .A3(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n721), .A3(new_n1020), .A4(new_n1018), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n725), .B1(new_n720), .B2(new_n724), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(new_n716), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n752), .A2(new_n763), .A3(new_n765), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1010), .B1(new_n1030), .B2(new_n767), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1008), .B(new_n1009), .C1(new_n1031), .C2(new_n771), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n231), .A2(new_n830), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n828), .C1(new_n212), .C2(new_n455), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n839), .B1(new_n1034), .B2(KEYINPUT110), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(KEYINPUT110), .B2(new_n1034), .ZN(new_n1036));
  INV_X1    g0836(.A(G283), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n513), .B1(new_n1037), .B2(new_n793), .C1(new_n808), .C2(new_n543), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n797), .A2(new_n626), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1039), .A2(KEYINPUT46), .B1(G107), .B2(new_n804), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(KEYINPUT46), .B2(new_n1039), .C1(new_n517), .C2(new_n788), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1038), .B(new_n1041), .C1(G317), .C2(new_n811), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n822), .A2(new_n617), .B1(new_n794), .B2(new_n800), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(KEYINPUT111), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT111), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n803), .A2(new_n316), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n851), .B2(new_n800), .C1(new_n788), .C2(new_n819), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n322), .B1(new_n793), .B2(new_n377), .C1(new_n234), .C2(new_n797), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G137), .B2(new_n811), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n365), .B2(new_n808), .C1(new_n850), .C2(new_n783), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1045), .A2(new_n1047), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n775), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n841), .B2(new_n1002), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1032), .A2(KEYINPUT112), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT112), .B1(new_n1032), .B2(new_n1057), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(G387));
  OAI21_X1  g0861(.A(KEYINPUT113), .B1(new_n1028), .B2(new_n729), .ZN(new_n1062));
  OAI21_X1  g0862(.A(KEYINPUT114), .B1(new_n767), .B2(new_n1026), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT113), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1027), .A2(new_n1064), .A3(new_n728), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT114), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1026), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n753), .C2(new_n766), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n730), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n836), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(G107), .B2(new_n212), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n228), .A2(G45), .ZN(new_n1073));
  AOI211_X1 g0873(.A(G45), .B(new_n1070), .C1(G68), .C2(G77), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n335), .A2(G50), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n831), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1072), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n772), .B1(new_n1078), .B2(new_n829), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n788), .A2(new_n335), .B1(new_n819), .B2(new_n800), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n797), .A2(new_n365), .B1(new_n793), .B2(new_n316), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1080), .A2(new_n513), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G97), .A2(new_n809), .B1(new_n811), .B2(G150), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n782), .A2(G50), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n454), .A2(new_n804), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n787), .A2(G311), .B1(new_n848), .B2(G303), .ZN(new_n1087));
  INV_X1    g0887(.A(G317), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(new_n784), .B2(new_n800), .C1(new_n822), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n797), .A2(new_n517), .B1(new_n803), .B2(new_n1037), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n268), .B1(new_n811), .B2(G326), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n626), .C2(new_n808), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n1098), .B2(new_n775), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n718), .A2(new_n719), .A3(new_n827), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n771), .B2(new_n1026), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1069), .A2(new_n1101), .ZN(G393));
  XNOR2_X1  g0902(.A(new_n1021), .B(new_n721), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1030), .B(new_n728), .C1(new_n1103), .C2(new_n1028), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n993), .A2(new_n827), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n240), .A2(new_n830), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n828), .C1(new_n543), .C2(new_n212), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n839), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n788), .A2(new_n377), .B1(new_n803), .B2(new_n365), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n268), .B1(new_n316), .B2(new_n797), .C1(new_n335), .C2(new_n793), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n859), .C1(new_n851), .C2(new_n810), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n782), .A2(G159), .B1(G150), .B2(new_n801), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n782), .A2(G311), .B1(G317), .B2(new_n801), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n788), .A2(new_n617), .B1(new_n803), .B2(new_n626), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n489), .B1(new_n793), .B2(new_n517), .C1(new_n1037), .C2(new_n797), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n444), .B2(new_n808), .C1(new_n784), .C2(new_n810), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1110), .B1(new_n1123), .B2(new_n775), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1103), .A2(new_n771), .B1(new_n1105), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1104), .A2(new_n1125), .ZN(G390));
  INV_X1    g0926(.A(new_n977), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n970), .B1(new_n1127), .B2(new_n978), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n950), .A2(new_n953), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n964), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT39), .B1(new_n1131), .B2(new_n968), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n937), .A2(new_n938), .A3(new_n962), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT106), .B1(new_n346), .B2(new_n300), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT37), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n931), .A2(new_n1136), .A3(new_n944), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(new_n930), .B1(new_n946), .B2(KEYINPUT107), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n359), .A2(new_n657), .A3(new_n361), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1139), .A2(new_n949), .B1(new_n951), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n968), .B1(new_n1141), .B2(KEYINPUT38), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n761), .A2(new_n710), .A3(new_n872), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n869), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n970), .B1(new_n1144), .B2(new_n978), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n751), .A2(G330), .A3(new_n874), .A4(new_n978), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1134), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n903), .A2(G330), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n899), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1128), .B1(new_n963), .B2(new_n969), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1148), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n479), .A2(new_n1150), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n985), .A2(new_n1157), .A3(new_n671), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n750), .B(new_n749), .C1(KEYINPUT94), .C2(new_n746), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n748), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n874), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n979), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1151), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1127), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n979), .B1(new_n1149), .B2(new_n873), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1147), .A2(new_n869), .A3(new_n1143), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1158), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n729), .B1(new_n1156), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1148), .A2(new_n1155), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1148), .A2(new_n1155), .A3(new_n771), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n825), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1173));
  INV_X1    g0973(.A(G137), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n788), .A2(new_n1174), .B1(new_n803), .B2(new_n819), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n783), .A2(new_n846), .B1(new_n377), .B2(new_n808), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n798), .A2(G150), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n1179), .B2(new_n800), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n811), .A2(G125), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n793), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n322), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1185));
  OR4_X1    g0985(.A1(new_n1175), .A2(new_n1176), .A3(new_n1180), .A4(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n788), .A2(new_n444), .B1(new_n803), .B2(new_n365), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G283), .B2(new_n801), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n489), .B1(new_n793), .B2(new_n543), .C1(new_n263), .C2(new_n797), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G68), .B2(new_n809), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n782), .A2(G116), .B1(G294), .B2(new_n811), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n776), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n839), .B(new_n1193), .C1(new_n335), .C2(new_n864), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1173), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1172), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(G378));
  AOI21_X1  g0998(.A(KEYINPUT40), .B1(new_n974), .B2(new_n904), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n955), .A2(G330), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n381), .A2(new_n912), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n395), .B(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1199), .A2(new_n1200), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n715), .B1(new_n1142), .B2(new_n942), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1208), .B2(new_n941), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n984), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1206), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n983), .A2(new_n973), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n941), .A3(new_n1205), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n971), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n985), .A2(new_n1157), .A3(new_n671), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT121), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1170), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1218), .A3(KEYINPUT57), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n728), .B(new_n1219), .C1(new_n1220), .C2(KEYINPUT57), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1206), .A2(new_n825), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n772), .B1(new_n865), .B2(G50), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G41), .B(new_n268), .C1(G77), .C2(new_n798), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT118), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n782), .A2(G107), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT119), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1049), .B1(new_n626), .B2(new_n800), .C1(new_n788), .C2(new_n543), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n809), .A2(G58), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n1037), .B2(new_n810), .C1(new_n455), .C2(new_n793), .ZN(new_n1230));
  OR4_X1    g1030(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT58), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n797), .A2(new_n1183), .B1(new_n793), .B2(new_n1174), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G132), .B2(new_n787), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n801), .A2(G125), .B1(new_n804), .B2(G150), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n783), .C2(new_n1179), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT59), .Z(new_n1239));
  NOR2_X1   g1039(.A1(G33), .A2(G41), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT117), .Z(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n811), .B2(G124), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n819), .B2(new_n808), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT120), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1241), .B(new_n377), .C1(new_n268), .C2(G41), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1233), .A2(new_n1234), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1223), .B1(new_n1247), .B2(new_n775), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1215), .A2(new_n771), .B1(new_n1222), .B2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1221), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT122), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1221), .A2(new_n1249), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(G375));
  NAND3_X1  g1056(.A1(new_n1164), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1258), .A2(new_n1010), .A3(new_n1167), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n771), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n772), .B1(new_n865), .B2(G68), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n822), .A2(new_n1174), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n788), .A2(new_n1183), .B1(new_n377), .B2(new_n803), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G132), .B2(new_n801), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n811), .A2(G128), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n797), .A2(new_n819), .B1(new_n793), .B2(new_n850), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n513), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1229), .A3(new_n1266), .A4(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n787), .A2(G116), .B1(new_n801), .B2(G294), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n322), .B1(new_n798), .B2(G97), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n444), .C2(new_n793), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n782), .A2(G283), .B1(G303), .B2(new_n811), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n1085), .C1(new_n365), .C2(new_n808), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1263), .A2(new_n1269), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1262), .B1(new_n1275), .B2(new_n775), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n978), .B2(new_n826), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1259), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT123), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(G381));
  AOI21_X1  g1081(.A(new_n1196), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1069), .A2(new_n843), .A3(new_n1101), .ZN(new_n1283));
  OR3_X1    g1083(.A1(G390), .A2(G384), .A3(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(G387), .A2(G381), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1255), .A2(new_n1282), .A3(new_n1285), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n1255), .A2(new_n1282), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n708), .A2(G213), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(KEYINPUT124), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G407), .B(G213), .C1(new_n1287), .C2(new_n1290), .ZN(G409));
  NOR3_X1   g1091(.A1(new_n1207), .A2(new_n1209), .A3(new_n984), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1211), .A2(new_n1213), .B1(new_n1212), .B2(new_n971), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT57), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1170), .A2(new_n1217), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n728), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1249), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(new_n1010), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1215), .A2(new_n771), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1222), .A2(new_n1248), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1282), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1290), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1260), .A2(new_n1216), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1257), .B1(new_n1167), .B2(new_n1308), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n728), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1278), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1307), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1312), .A2(new_n1314), .A3(new_n1307), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(G2897), .A3(new_n1289), .A4(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1289), .A2(G2897), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1317), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1315), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1320), .A2(new_n1315), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1306), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1069), .A2(new_n843), .A3(new_n1101), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n843), .B1(new_n1069), .B2(new_n1101), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1327), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G393), .A2(G396), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(KEYINPUT126), .A3(new_n1283), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1032), .A2(new_n1057), .A3(G390), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G390), .B1(new_n1032), .B2(new_n1057), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1334), .A2(new_n1336), .A3(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1330), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1335), .B1(new_n1340), .B2(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G390), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1342));
  AOI22_X1  g1142(.A1(new_n1339), .A2(new_n1341), .B1(G387), .B2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1289), .B1(new_n1298), .B2(new_n1304), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1325), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1323), .A2(new_n1326), .A3(new_n1343), .A4(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT62), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1344), .A2(new_n1348), .A3(new_n1345), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1350), .B1(new_n1344), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1348), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1349), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1347), .B1(new_n1354), .B2(new_n1343), .ZN(G405));
  NOR2_X1   g1155(.A1(new_n1250), .A2(new_n1282), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1339), .A2(new_n1341), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1060), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1342), .A2(new_n1359), .A3(new_n1058), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1358), .A2(new_n1360), .A3(new_n1325), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1325), .B1(new_n1358), .B2(new_n1360), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1287), .B(new_n1357), .C1(new_n1361), .C2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1336), .B1(new_n1334), .B2(new_n1338), .ZN(new_n1364));
  NOR3_X1   g1164(.A1(new_n1340), .A2(new_n1337), .A3(new_n1335), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1360), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1345), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1343), .A2(new_n1325), .ZN(new_n1368));
  AOI21_X1  g1168(.A(G378), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n1367), .B(new_n1368), .C1(new_n1369), .C2(new_n1356), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1363), .A2(new_n1370), .ZN(G402));
endmodule


