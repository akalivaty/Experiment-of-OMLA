//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n204), .A2(G50), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT67), .B(G238), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n203), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G107), .A2(G264), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n213), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n216), .B1(new_n222), .B2(new_n223), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT66), .B(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(new_n254), .B2(new_n255), .C1(new_n205), .C2(new_n211), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(G50), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n210), .B2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n263), .A2(new_n265), .B1(new_n264), .B2(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n273), .A3(G274), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT69), .Z(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G223), .A3(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G77), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n273), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n279), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n268), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(G190), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT10), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(new_n279), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n302), .A3(new_n309), .A4(new_n268), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n307), .A2(new_n312), .B1(new_n260), .B2(new_n266), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n299), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G244), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n274), .B1(new_n317), .B2(new_n277), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n289), .A2(G1698), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n319), .B1(new_n320), .B2(new_n289), .C1(new_n321), .C2(new_n224), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n258), .B1(G33), .B2(G41), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n324), .A2(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n206), .B1(new_n210), .B2(G20), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n263), .A2(new_n326), .B1(new_n206), .B2(new_n262), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT72), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n254), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n255), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n251), .B1(new_n220), .B2(G77), .ZN(new_n332));
  INV_X1    g0132(.A(new_n329), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT72), .A3(G33), .A4(new_n253), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n259), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n327), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n324), .B2(G169), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n324), .B2(G190), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n300), .B2(new_n324), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n311), .A2(new_n316), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n283), .A2(new_n288), .A3(G232), .A4(G1698), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n283), .A2(new_n288), .A3(G226), .A4(new_n290), .ZN(new_n346));
  INV_X1    g0146(.A(G97), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT73), .B1(new_n285), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(G33), .A3(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n323), .ZN(new_n353));
  INV_X1    g0153(.A(new_n274), .ZN(new_n354));
  INV_X1    g0154(.A(G238), .ZN(new_n355));
  INV_X1    g0155(.A(new_n277), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n277), .A2(KEYINPUT74), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n353), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(G190), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n253), .A2(G33), .A3(G77), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n203), .A2(G20), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT76), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n211), .A2(new_n285), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n264), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT76), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n259), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT11), .B(new_n259), .C1(new_n370), .C2(new_n371), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT12), .B1(new_n261), .B2(G68), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n203), .B1(new_n210), .B2(G20), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n376), .A2(new_n377), .B1(new_n263), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n365), .A2(new_n374), .A3(new_n375), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n362), .A2(new_n364), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n300), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n362), .A2(new_n364), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT75), .A3(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n374), .A2(new_n375), .A3(new_n379), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT14), .B1(new_n382), .B2(new_n312), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n362), .A2(G179), .A3(new_n364), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n255), .B1(new_n210), .B2(G20), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n263), .B1(new_n262), .B2(new_n255), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n281), .A2(new_n282), .A3(G20), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n281), .A2(new_n282), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n400), .A2(new_n253), .A3(new_n398), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT77), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n286), .A2(new_n211), .A3(new_n287), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n203), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT77), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n253), .A3(new_n398), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G58), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n211), .B1(new_n204), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n251), .A2(G159), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT78), .A3(new_n412), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n336), .B1(new_n408), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n398), .A2(new_n211), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n283), .B2(new_n288), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n398), .B1(new_n400), .B2(new_n253), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(new_n203), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n412), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n396), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT80), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n275), .A2(G1698), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n431), .B1(G223), .B2(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n323), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n274), .B1(new_n235), .B2(new_n277), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n300), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n273), .B1(new_n432), .B2(new_n433), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n439), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n429), .A2(KEYINPUT80), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n428), .A2(new_n430), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n419), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n427), .A3(new_n259), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n442), .A3(new_n395), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT80), .A3(new_n429), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n395), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n312), .B1(new_n435), .B2(new_n437), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n439), .A2(new_n436), .A3(new_n314), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  AOI211_X1 g0258(.A(KEYINPUT18), .B(new_n456), .C1(new_n448), .C2(new_n395), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT79), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT18), .B1(new_n428), .B2(new_n456), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n453), .A2(new_n452), .A3(new_n457), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n451), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n344), .A2(new_n393), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n262), .A2(new_n347), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n210), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n261), .A2(new_n469), .A3(new_n258), .A4(new_n257), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(new_n347), .ZN(new_n471));
  AND2_X1   g0271(.A1(G97), .A2(G107), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(KEYINPUT6), .B2(new_n347), .ZN(new_n476));
  XNOR2_X1  g0276(.A(G97), .B(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT82), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n474), .B(new_n480), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n220), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n424), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(G107), .C1(new_n289), .C2(new_n422), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n251), .A2(G77), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n471), .B1(new_n486), .B2(new_n259), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n283), .A2(new_n288), .A3(G250), .A4(G1698), .ZN(new_n488));
  AND2_X1   g0288(.A1(KEYINPUT4), .A2(G244), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n283), .A2(new_n288), .A3(new_n290), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(new_n290), .C1(new_n281), .C2(new_n282), .ZN(new_n492));
  XOR2_X1   g0292(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n323), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n210), .B(G45), .C1(new_n269), .C2(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(KEYINPUT84), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n270), .A2(G1), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G257), .B(new_n273), .C1(new_n499), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n500), .A3(new_n503), .ZN(new_n507));
  INV_X1    g0307(.A(G274), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n221), .B2(new_n272), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n497), .A4(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n496), .A2(new_n511), .A3(G190), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n496), .A2(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(G200), .ZN(new_n515));
  AOI211_X1 g0315(.A(KEYINPUT85), .B(new_n300), .C1(new_n496), .C2(new_n511), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n487), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n486), .A2(new_n259), .ZN(new_n518));
  INV_X1    g0318(.A(new_n471), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n496), .A2(new_n511), .A3(new_n314), .ZN(new_n521));
  AOI21_X1  g0321(.A(G169), .B1(new_n496), .B2(new_n511), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n286), .A2(new_n287), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n317), .A2(G1698), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(G238), .C2(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n285), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n273), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n273), .A2(G274), .A3(new_n501), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n509), .A2(new_n535), .A3(new_n501), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(G250), .B1(new_n270), .B2(G1), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n221), .B2(new_n272), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT87), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT87), .ZN(new_n542));
  AOI211_X1 g0342(.A(new_n542), .B(new_n539), .C1(new_n534), .C2(new_n536), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n314), .B(new_n532), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n470), .A2(new_n329), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT88), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n217), .A2(new_n219), .A3(G33), .A4(G97), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n525), .A2(new_n253), .A3(G68), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT19), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n253), .B1(new_n553), .B2(new_n473), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n259), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n329), .A2(new_n262), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n546), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n535), .B1(new_n509), .B2(new_n501), .ZN(new_n558));
  AND4_X1   g0358(.A1(new_n535), .A2(new_n273), .A3(G274), .A4(new_n501), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n540), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n542), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n537), .A2(KEYINPUT87), .A3(new_n540), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n531), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n544), .B(new_n557), .C1(new_n563), .C2(G169), .ZN(new_n564));
  OAI211_X1 g0364(.A(G190), .B(new_n532), .C1(new_n541), .C2(new_n543), .ZN(new_n565));
  OR2_X1    g0365(.A1(new_n470), .A2(new_n553), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n555), .A2(new_n556), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n567), .C1(new_n563), .C2(new_n300), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n517), .A2(new_n524), .A3(new_n564), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n283), .B2(new_n288), .ZN(new_n571));
  INV_X1    g0371(.A(G264), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G1698), .ZN(new_n573));
  OAI221_X1 g0373(.A(new_n573), .B1(G257), .B2(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n323), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G270), .B(new_n273), .C1(new_n499), .C2(new_n504), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n510), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n262), .A2(new_n528), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n470), .B2(new_n528), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n285), .A2(G97), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n253), .A2(new_n491), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n257), .A2(new_n258), .B1(G20), .B2(new_n528), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n578), .A2(new_n588), .A3(new_n314), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n312), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(new_n578), .ZN(new_n592));
  INV_X1    g0392(.A(new_n580), .ZN(new_n593));
  INV_X1    g0393(.A(new_n587), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n582), .B2(new_n583), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n578), .A2(new_n596), .A3(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT21), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n589), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT22), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n293), .B2(new_n553), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n220), .A2(new_n603), .B1(KEYINPUT23), .B2(G107), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n525), .A2(new_n253), .A3(KEYINPUT22), .A4(G87), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n211), .B1(new_n529), .B2(KEYINPUT23), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT24), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n607), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n601), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n259), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n320), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT25), .B1(new_n262), .B2(new_n320), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n320), .B2(new_n470), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G264), .B(new_n273), .C1(new_n499), .C2(new_n504), .ZN(new_n619));
  INV_X1    g0419(.A(G257), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G1698), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G250), .B2(G1698), .ZN(new_n622));
  INV_X1    g0422(.A(G294), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n400), .B1(new_n285), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n323), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n510), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(new_n440), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(G200), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n613), .A2(new_n618), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(G169), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n314), .B2(new_n626), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n336), .B1(new_n608), .B2(new_n611), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n617), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n596), .B1(new_n578), .B2(G200), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n440), .B2(new_n578), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n599), .A2(new_n629), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n467), .A2(new_n569), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n316), .ZN(new_n638));
  INV_X1    g0438(.A(new_n311), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n391), .A2(new_n389), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n390), .B1(new_n384), .B2(G169), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n387), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n386), .B2(new_n340), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n444), .A2(new_n450), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n458), .A2(new_n459), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(KEYINPUT90), .A3(new_n646), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n638), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n517), .A2(new_n524), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n627), .A2(new_n628), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n653), .A2(new_n632), .A3(new_n617), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n599), .B2(new_n633), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n564), .A2(new_n568), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n656), .B2(new_n524), .ZN(new_n660));
  INV_X1    g0460(.A(new_n521), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n487), .A2(new_n661), .A3(new_n522), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n564), .A4(new_n568), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT89), .B1(new_n664), .B2(new_n564), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  INV_X1    g0466(.A(new_n564), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n666), .B(new_n667), .C1(new_n660), .C2(new_n663), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n658), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n651), .B1(new_n467), .B2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(new_n599), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n253), .A2(new_n210), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n588), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n592), .A2(new_n598), .ZN(new_n680));
  INV_X1    g0480(.A(new_n589), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n635), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT91), .Z(new_n685));
  INV_X1    g0485(.A(new_n633), .ZN(new_n686));
  INV_X1    g0486(.A(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n632), .B2(new_n617), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n629), .A2(new_n633), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n685), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n599), .A2(new_n687), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n686), .A2(new_n677), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n214), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G1), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n473), .A2(new_n553), .A3(new_n528), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n710), .B1(new_n223), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n667), .B1(new_n660), .B2(new_n663), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n687), .B1(new_n658), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n664), .A2(new_n564), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n666), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n687), .B1(new_n719), .B2(new_n658), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n715), .B1(new_n720), .B2(KEYINPUT29), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n569), .A2(new_n636), .A3(new_n687), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  AND4_X1   g0524(.A1(G179), .A2(new_n510), .A3(new_n619), .A4(new_n625), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n576), .A2(new_n577), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n496), .A4(new_n511), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n532), .B1(new_n541), .B2(new_n543), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n724), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT95), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n578), .A2(new_n314), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n563), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n728), .A2(KEYINPUT95), .A3(new_n314), .A4(new_n578), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n514), .A4(new_n626), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n687), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n723), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n722), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n721), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n712), .B1(new_n745), .B2(G1), .ZN(G364));
  AND2_X1   g0546(.A1(new_n253), .A2(G13), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n709), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n258), .B1(G20), .B2(new_n312), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n706), .A2(new_n293), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G355), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n214), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n706), .A2(new_n525), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n223), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n270), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n249), .A2(G45), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n253), .A2(new_n314), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(new_n440), .A3(new_n300), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G326), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n211), .A2(new_n440), .A3(new_n300), .A4(G179), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n289), .B1(G303), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n440), .A2(G200), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n253), .B1(new_n314), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n769), .B(new_n771), .C1(new_n623), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n767), .A2(G190), .A3(new_n300), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n766), .A2(new_n772), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G190), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n220), .A2(new_n300), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n779), .A2(G322), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n220), .A2(G200), .A3(new_n780), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n766), .A2(new_n440), .A3(new_n300), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n786), .B1(new_n793), .B2(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n773), .A2(new_n347), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n768), .B1(new_n775), .B2(G68), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n293), .B1(G87), .B2(new_n770), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n785), .A2(new_n320), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n779), .B2(G58), .ZN(new_n800));
  AND4_X1   g0600(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT32), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n781), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n782), .A2(KEYINPUT32), .A3(G159), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n793), .A2(G77), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n777), .A2(new_n794), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n754), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n750), .B1(new_n756), .B2(new_n765), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  INV_X1    g0610(.A(new_n753), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n683), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT98), .ZN(new_n813));
  INV_X1    g0613(.A(new_n750), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n685), .B(new_n814), .C1(G330), .C2(new_n683), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n340), .A2(new_n687), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n687), .A2(new_n337), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n339), .B1(new_n342), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n720), .B(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(new_n743), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n750), .B1(new_n821), .B2(new_n743), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n754), .A2(new_n751), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  INV_X1    g0626(.A(new_n785), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G87), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n623), .B2(new_n778), .C1(new_n829), .C2(new_n781), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n289), .B(new_n795), .C1(G107), .C2(new_n770), .ZN(new_n831));
  INV_X1    g0631(.A(new_n775), .ZN(new_n832));
  INV_X1    g0632(.A(new_n768), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n784), .B2(new_n832), .C1(new_n570), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n830), .B(new_n834), .C1(G116), .C2(new_n793), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n768), .A2(G137), .B1(G143), .B2(new_n779), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n832), .C1(new_n792), .C2(new_n803), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n773), .A2(new_n202), .ZN(new_n840));
  INV_X1    g0640(.A(new_n770), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n525), .B1(new_n785), .B2(new_n203), .C1(new_n841), .C2(new_n264), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G132), .C2(new_n782), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n835), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n750), .B1(G77), .B2(new_n826), .C1(new_n844), .C2(new_n808), .ZN(new_n845));
  INV_X1    g0645(.A(new_n820), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n751), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT100), .Z(new_n848));
  NOR2_X1   g0648(.A1(new_n824), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n479), .A2(new_n481), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT35), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n528), .B(new_n222), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(new_n852), .B2(new_n851), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT36), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n223), .A2(new_n206), .A3(new_n415), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(KEYINPUT102), .ZN(new_n860));
  INV_X1    g0660(.A(new_n201), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n859), .A2(KEYINPUT102), .B1(G68), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n210), .B(G13), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n414), .B(new_n418), .C1(new_n445), .C2(new_n446), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n421), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n396), .B1(new_n866), .B2(new_n420), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n449), .B1(new_n867), .B2(new_n456), .ZN(new_n868));
  INV_X1    g0668(.A(new_n676), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n453), .A2(new_n457), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n453), .A2(new_n676), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n449), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n870), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n465), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT38), .B(new_n876), .C1(new_n465), .C2(new_n877), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(KEYINPUT103), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n883), .A3(new_n879), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n872), .A2(new_n873), .A3(new_n449), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT104), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n875), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n888), .B2(new_n875), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n873), .B1(new_n644), .B2(new_n646), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n881), .B(new_n886), .C1(new_n894), .C2(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n392), .A2(new_n387), .A3(new_n677), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n646), .A2(new_n676), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n882), .A2(new_n884), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n387), .B(new_n687), .C1(new_n386), .C2(new_n392), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n387), .B1(new_n382), .B2(G190), .ZN(new_n903));
  INV_X1    g0703(.A(new_n385), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT75), .B1(new_n384), .B2(G200), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n387), .A2(new_n687), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n642), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n669), .A2(new_n677), .A3(new_n820), .ZN(new_n911));
  INV_X1    g0711(.A(new_n817), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n900), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n899), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n466), .B(new_n715), .C1(new_n720), .C2(KEYINPUT29), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n651), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n738), .A2(new_n687), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT31), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n629), .A2(new_n633), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n682), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(new_n652), .A3(new_n657), .A4(new_n677), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n924), .A3(new_n741), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n925), .A2(new_n909), .A3(new_n820), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n882), .A2(new_n926), .A3(new_n884), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n892), .A2(new_n893), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n890), .ZN(new_n931));
  INV_X1    g0731(.A(new_n881), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT106), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n881), .C1(new_n894), .C2(KEYINPUT38), .ZN(new_n935));
  AND4_X1   g0735(.A1(KEYINPUT40), .A2(new_n925), .A3(new_n820), .A4(new_n909), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n466), .A2(new_n925), .ZN(new_n939));
  OAI21_X1  g0739(.A(G330), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n918), .A2(new_n941), .B1(new_n210), .B2(new_n747), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n918), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n864), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OR2_X1    g0744(.A1(new_n567), .A2(new_n677), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n657), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n564), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n652), .B1(new_n487), .B2(new_n677), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n662), .A2(new_n687), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT42), .B1(new_n702), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n524), .B1(new_n949), .B2(new_n633), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n677), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n702), .A2(KEYINPUT42), .A3(new_n952), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n700), .A3(new_n951), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(new_n700), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n952), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n707), .B(new_n966), .Z(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n704), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT44), .B1(new_n704), .B2(new_n952), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n702), .A2(new_n703), .A3(new_n951), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT45), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n975), .A3(new_n964), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n700), .B1(new_n971), .B2(new_n974), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n698), .A2(KEYINPUT108), .A3(new_n701), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT108), .B1(new_n698), .B2(new_n701), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n685), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n685), .A3(new_n981), .A4(new_n982), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n976), .A2(new_n977), .A3(new_n987), .A4(new_n745), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n968), .B1(new_n988), .B2(new_n745), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n749), .A2(new_n210), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n962), .B(new_n965), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n755), .B1(new_n214), .B2(new_n329), .C1(new_n761), .C2(new_n241), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(new_n750), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n841), .A2(new_n995), .A3(new_n528), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT46), .B1(new_n770), .B2(G116), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n996), .A2(new_n525), .A3(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n832), .B2(new_n623), .C1(new_n829), .C2(new_n833), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n792), .A2(new_n784), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n773), .A2(new_n320), .B1(new_n781), .B2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n778), .A2(new_n570), .B1(new_n347), .B2(new_n785), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n773), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(G68), .ZN(new_n1006));
  INV_X1    g0806(.A(G137), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n781), .C1(new_n778), .C2(new_n837), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n775), .A2(G159), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n768), .A2(G143), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n827), .A2(G77), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n293), .B1(G58), .B2(new_n770), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1008), .B(new_n1013), .C1(new_n201), .C2(new_n793), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1004), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n994), .B1(new_n811), .B2(new_n947), .C1(new_n1016), .C2(new_n808), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n992), .A2(new_n1017), .ZN(G387));
  NOR2_X1   g0818(.A1(new_n987), .A2(new_n745), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n987), .A2(new_n745), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n707), .A3(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n238), .A2(new_n270), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(new_n760), .B1(new_n710), .B2(new_n757), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n331), .B2(new_n264), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n270), .B1(new_n203), .B2(new_n206), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n710), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1024), .A2(new_n1029), .B1(G107), .B2(new_n214), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n814), .B1(new_n1030), .B2(new_n755), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1005), .A2(new_n333), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n837), .B2(new_n781), .C1(new_n778), .C2(new_n264), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n525), .B1(new_n841), .B2(new_n206), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G97), .B2(new_n827), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n832), .B2(new_n255), .C1(new_n803), .C2(new_n833), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(G68), .C2(new_n793), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n775), .A2(G311), .B1(G317), .B2(new_n779), .ZN(new_n1038));
  INV_X1    g0838(.A(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n833), .C1(new_n792), .C2(new_n570), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1005), .A2(G283), .B1(new_n770), .B2(G294), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n525), .B1(new_n782), .B2(G326), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n528), .B2(new_n785), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1046), .B2(KEYINPUT49), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1037), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1031), .B1(new_n1051), .B2(new_n808), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n699), .B2(new_n753), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n987), .B2(new_n991), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1022), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT110), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1021), .A2(new_n707), .ZN(new_n1058));
  OAI211_X1 g0858(.A(KEYINPUT110), .B(new_n1054), .C1(new_n1058), .C2(new_n1019), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(G393));
  NAND3_X1  g0860(.A1(new_n976), .A2(new_n991), .A3(new_n977), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n246), .A2(new_n761), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n755), .B1(new_n347), .B2(new_n214), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n832), .A2(new_n570), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n289), .B(new_n799), .C1(G283), .C2(new_n770), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n528), .B2(new_n773), .C1(new_n1039), .C2(new_n781), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G294), .C2(new_n793), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n768), .A2(G317), .B1(G311), .B2(new_n779), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n768), .A2(G150), .B1(G159), .B2(new_n779), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n1005), .A2(G77), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n400), .B1(new_n770), .B2(G68), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n782), .A2(G143), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1072), .A2(new_n828), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n832), .A2(new_n861), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n793), .C2(new_n331), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1067), .A2(new_n1069), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n750), .B1(new_n1062), .B2(new_n1063), .C1(new_n1078), .C2(new_n808), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT111), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n811), .B2(new_n951), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT112), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT112), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1061), .A2(new_n1084), .A3(new_n1081), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n988), .A2(new_n707), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n976), .A2(new_n977), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1021), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1086), .A2(new_n1090), .ZN(G390));
  NAND3_X1  g0891(.A1(new_n902), .A2(KEYINPUT113), .A3(new_n908), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n642), .A2(new_n906), .A3(new_n907), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n907), .B1(new_n642), .B2(new_n906), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n819), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n714), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1092), .B(new_n1096), .C1(new_n1098), .C2(new_n817), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1099), .A2(new_n933), .A3(new_n897), .A4(new_n935), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n911), .A2(new_n912), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n898), .B1(new_n1101), .B2(new_n909), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n896), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n925), .A2(new_n909), .A3(new_n820), .A4(G330), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1100), .C1(new_n1102), .C2(new_n896), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n991), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n750), .B1(new_n826), .B2(new_n331), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT117), .Z(new_n1110));
  AOI22_X1  g0910(.A1(G107), .A2(new_n775), .B1(new_n768), .B2(G283), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n792), .B2(new_n347), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT119), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n293), .B1(new_n785), .B2(new_n203), .C1(new_n841), .C2(new_n553), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1072), .B1(new_n623), .B2(new_n781), .C1(new_n778), .C2(new_n528), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  AOI21_X1  g0917(.A(new_n293), .B1(new_n827), .B2(new_n201), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n793), .A2(new_n1117), .B1(KEYINPUT118), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(KEYINPUT118), .B2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n770), .A2(G150), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT53), .Z(new_n1122));
  AOI22_X1  g0922(.A1(new_n779), .A2(G132), .B1(new_n782), .B2(G125), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n803), .C2(new_n773), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n768), .A2(G128), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n832), .B2(new_n1007), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1116), .A2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1110), .B1(new_n808), .B2(new_n1128), .C1(new_n896), .C2(new_n752), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1108), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT120), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n466), .A2(new_n742), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n916), .A2(new_n651), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n742), .A2(new_n820), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n817), .B1(new_n714), .B2(new_n1097), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1104), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1096), .A2(new_n1092), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n925), .A2(G330), .A3(new_n820), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT114), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n1104), .A4(new_n1136), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n909), .B1(new_n742), .B2(new_n820), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1101), .B1(new_n1145), .B2(new_n1105), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1134), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1106), .A2(new_n1147), .A3(new_n1107), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n707), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(KEYINPUT115), .A3(new_n707), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1151), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1132), .A2(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(new_n1134), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n929), .A2(new_n937), .A3(G330), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n915), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n267), .A2(new_n676), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n311), .A2(new_n316), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n311), .B2(new_n316), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1168), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT122), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n899), .B(new_n914), .C1(new_n938), .C2(new_n722), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1164), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1173), .B1(new_n1164), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1162), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n708), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1162), .B(KEYINPUT57), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT123), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1164), .A2(new_n1174), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1172), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1164), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT123), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT57), .A4(new_n1162), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1179), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1171), .A2(new_n751), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n750), .B1(new_n826), .B2(new_n201), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n827), .A2(G58), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n320), .B2(new_n778), .C1(new_n784), .C2(new_n781), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n400), .A2(new_n269), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G77), .B2(new_n770), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1006), .A2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n832), .B2(new_n347), .C1(new_n528), .C2(new_n833), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1192), .B(new_n1196), .C1(new_n333), .C2(new_n793), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT58), .Z(new_n1198));
  OAI211_X1 g0998(.A(new_n1193), .B(new_n264), .C1(G33), .C2(G41), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G125), .A2(new_n768), .B1(new_n775), .B2(G132), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n779), .A2(G128), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1005), .A2(G150), .B1(new_n770), .B2(new_n1117), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G137), .B2(new_n793), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n285), .B(new_n269), .C1(new_n785), .C2(new_n803), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G124), .B2(new_n782), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1198), .B(new_n1199), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT121), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n808), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1190), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1185), .A2(new_n991), .B1(new_n1189), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1188), .A2(new_n1216), .ZN(G375));
  OAI21_X1  g1017(.A(new_n750), .B1(new_n826), .B2(G68), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n289), .B1(G97), .B2(new_n770), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1011), .B(new_n1219), .C1(new_n832), .C2(new_n528), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G294), .B2(new_n768), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1032), .B1(new_n570), .B2(new_n781), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G283), .B2(new_n779), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(new_n320), .C2(new_n792), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n768), .A2(G132), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n775), .A2(new_n1117), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n400), .B1(new_n770), .B2(G159), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1191), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n779), .A2(G137), .B1(new_n782), .B2(G128), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n264), .B2(new_n773), .C1(new_n792), .C2(new_n837), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1224), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT125), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n808), .B1(new_n1231), .B2(KEYINPUT125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1218), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1139), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n752), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n990), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1134), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT124), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1153), .A2(new_n967), .A3(new_n1156), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1239), .B1(new_n1243), .B2(new_n1244), .ZN(G381));
  AOI22_X1  g1045(.A1(new_n1083), .A2(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n849), .ZN(new_n1247));
  INV_X1    g1047(.A(G396), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1057), .A2(new_n1248), .A3(new_n1059), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1247), .A2(new_n1249), .A3(G387), .A4(G381), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1132), .A2(new_n1159), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1216), .A4(new_n1188), .ZN(G407));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G343), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G375), .C2(new_n1255), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n1188), .A2(G378), .A3(new_n1216), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1216), .B1(new_n968), .B2(new_n1177), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT126), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1254), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1241), .A2(new_n1242), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1240), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n708), .B1(new_n1265), .B2(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G384), .A3(new_n1239), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1267), .B2(new_n1239), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1257), .A2(new_n1259), .A3(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1261), .A2(new_n1262), .A3(new_n1271), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n1262), .A3(new_n1273), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1270), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1278), .A2(new_n1268), .A3(G2897), .A4(new_n1254), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1254), .A2(G2897), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1246), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT127), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT110), .B1(new_n1022), .B2(new_n1054), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1059), .ZN(new_n1287));
  OAI21_X1  g1087(.A(G396), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1249), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G390), .A2(new_n992), .A3(new_n1017), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1285), .A2(new_n1289), .B1(new_n1290), .B2(new_n1284), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  AND4_X1   g1092(.A1(new_n1292), .A2(new_n1289), .A3(new_n1284), .A4(new_n1290), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(KEYINPUT61), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1254), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1276), .A2(new_n1283), .A3(new_n1295), .A4(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1296), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1274), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1296), .A2(KEYINPUT62), .A3(new_n1271), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1301), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1294), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1298), .B1(new_n1305), .B2(new_n1306), .ZN(G405));
  XNOR2_X1  g1107(.A(G375), .B(G378), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1271), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1310), .A2(new_n1294), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1294), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


