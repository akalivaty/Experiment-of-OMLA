//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(KEYINPUT0), .B2(new_n213), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n233));
  INV_X1    g0033(.A(G226), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n233), .B1(new_n202), .B2(new_n234), .ZN(new_n235));
  NOR4_X1   g0035(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  OR2_X1    g0036(.A1(new_n236), .A2(new_n208), .ZN(new_n237));
  AND2_X1   g0037(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n239));
  NOR3_X1   g0039(.A1(new_n221), .A2(new_n238), .A3(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G68), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n254), .B(new_n255), .Z(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  NAND2_X1  g0057(.A1(new_n208), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n214), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n209), .A2(new_n207), .A3(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n261), .A2(new_n262), .B1(new_n202), .B2(new_n260), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n208), .B2(G33), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n207), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(G20), .B2(new_n203), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n263), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT72), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n282), .B1(new_n283), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n264), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n264), .B2(new_n287), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(new_n294), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(G226), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n275), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(KEYINPUT72), .A3(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G190), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n274), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(new_n273), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n300), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n310), .A2(new_n311), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n297), .A2(G244), .ZN(new_n317));
  INV_X1    g0117(.A(new_n280), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G107), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n280), .A2(G232), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n319), .B1(new_n284), .B2(new_n230), .C1(G1698), .C2(new_n320), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n296), .B(new_n317), .C1(new_n321), .C2(new_n289), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  INV_X1    g0123(.A(new_n266), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT15), .B(G87), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n325), .A2(new_n326), .B1(new_n267), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n259), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n283), .B1(new_n206), .B2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n261), .A2(new_n331), .B1(new_n283), .B2(new_n260), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n322), .A2(new_n312), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n322), .A2(G190), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n333), .C1(new_n301), .C2(new_n322), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n306), .A2(new_n316), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n316), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(new_n320), .C2(new_n281), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n289), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n296), .B1(G238), .B2(new_n297), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G169), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n354), .A2(G179), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n358), .A3(G169), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n260), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G68), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n363), .A2(KEYINPUT75), .A3(KEYINPUT12), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT75), .B1(new_n363), .B2(KEYINPUT12), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(KEYINPUT12), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n206), .A2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n261), .A2(G68), .A3(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n231), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n283), .B2(new_n267), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n259), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT11), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n350), .B2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n342), .A2(new_n343), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT76), .B(G33), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n278), .B1(new_n382), .B2(new_n276), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G223), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n234), .B2(G1698), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n385), .B1(G33), .B2(G87), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n288), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n297), .A2(G232), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n295), .ZN(new_n389));
  OAI21_X1  g0189(.A(G169), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n296), .B1(G232), .B2(new_n297), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(G179), .C1(new_n288), .C2(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G58), .A2(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n207), .B1(new_n216), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(G159), .B2(new_n269), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n207), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n383), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n277), .A2(KEYINPUT76), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G33), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n276), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n278), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT77), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n278), .C1(new_n382), .C2(new_n276), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n207), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n400), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n397), .C1(new_n411), .C2(new_n231), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n279), .A2(new_n207), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n410), .B(new_n413), .C1(new_n382), .C2(new_n276), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n405), .A2(new_n413), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n398), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n397), .B1(new_n417), .B2(new_n231), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n420), .A3(new_n259), .ZN(new_n421));
  INV_X1    g0221(.A(new_n261), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n324), .A2(new_n368), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n422), .A2(new_n423), .B1(new_n361), .B2(new_n324), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n394), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT18), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n391), .B1(new_n386), .B2(new_n288), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n301), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G190), .B2(new_n428), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n381), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT82), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT81), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n383), .A2(new_n440), .A3(G244), .A4(new_n281), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT4), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G244), .B(new_n281), .C1(new_n404), .C2(new_n405), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT81), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n435), .B1(new_n446), .B2(new_n288), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n442), .A3(new_n441), .ZN(new_n448));
  INV_X1    g0248(.A(new_n439), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n288), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n206), .B(G45), .C1(new_n452), .C2(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(KEYINPUT83), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n289), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G257), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT84), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n460), .A3(new_n292), .A4(new_n457), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n457), .A2(new_n467), .A3(new_n292), .A4(new_n453), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n470), .A3(new_n312), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n447), .A2(new_n451), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n448), .A2(new_n449), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n289), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n459), .A2(new_n470), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n307), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G97), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT80), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  AOI22_X1  g0283(.A1(KEYINPUT79), .A2(new_n483), .B1(new_n225), .B2(G107), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(KEYINPUT79), .B2(new_n483), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n482), .B(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n417), .A2(new_n480), .B1(new_n283), .B2(new_n270), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n259), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n361), .A2(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n206), .A2(G33), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n265), .A2(new_n361), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n473), .A2(new_n479), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT85), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n473), .A2(new_n479), .A3(KEYINPUT85), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n494), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n435), .B(new_n288), .C1(new_n448), .C2(new_n449), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n501), .A2(new_n502), .A3(new_n476), .ZN(new_n503));
  OAI221_X1 g0303(.A(new_n500), .B1(new_n378), .B2(new_n478), .C1(new_n503), .C2(new_n301), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n226), .A2(G1698), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G250), .B2(G1698), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n402), .A2(G33), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n277), .A2(KEYINPUT76), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT3), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n278), .ZN(new_n511));
  INV_X1    g0311(.A(G294), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n382), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n289), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n518));
  OAI211_X1 g0318(.A(G264), .B(new_n288), .C1(new_n455), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n457), .A2(new_n453), .A3(new_n467), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT90), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(G264), .A4(new_n288), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n517), .A2(new_n524), .A3(new_n312), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n401), .A2(new_n403), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n405), .B1(new_n526), .B2(KEYINPUT3), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n527), .A2(new_n507), .B1(new_n512), .B2(new_n382), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n461), .A2(new_n469), .B1(new_n528), .B2(new_n289), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n307), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT91), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n207), .B(G87), .C1(new_n404), .C2(new_n405), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n223), .A2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n280), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT23), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n207), .B2(G107), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n480), .A2(KEYINPUT23), .A3(G20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n526), .A2(G116), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(G20), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n532), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n537), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n533), .B2(KEYINPUT22), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n548), .A2(KEYINPUT24), .A3(new_n544), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n259), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT25), .B1(new_n260), .B2(new_n480), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n480), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n492), .A2(G107), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n514), .B(new_n519), .C1(new_n515), .C2(new_n516), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G169), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT91), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n520), .A2(new_n523), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n529), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n558), .C1(new_n560), .C2(new_n312), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n531), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT92), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n531), .A2(new_n555), .A3(new_n561), .A4(KEYINPUT92), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n550), .A2(new_n554), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n517), .A2(new_n524), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n568), .A2(G200), .B1(G190), .B2(new_n556), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(KEYINPUT93), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT93), .ZN(new_n571));
  INV_X1    g0371(.A(new_n556), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n301), .A2(new_n560), .B1(new_n572), .B2(new_n378), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n555), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n463), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n224), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n288), .C1(G274), .C2(new_n577), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G244), .B(G1698), .C1(new_n404), .C2(new_n405), .ZN(new_n581));
  OAI211_X1 g0381(.A(G238), .B(new_n281), .C1(new_n404), .C2(new_n405), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n543), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n583), .B2(new_n289), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n584), .A2(G169), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n312), .ZN(new_n586));
  INV_X1    g0386(.A(new_n327), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n361), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n492), .A2(new_n587), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n383), .A2(new_n207), .A3(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n207), .B1(new_n345), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n223), .A2(new_n225), .A3(new_n480), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n593), .A2(new_n594), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n589), .B(new_n590), .C1(new_n597), .C2(new_n265), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n585), .A2(new_n586), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n584), .A2(G190), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n265), .B1(new_n591), .B2(new_n596), .ZN(new_n602));
  AND4_X1   g0402(.A1(G87), .A2(new_n265), .A3(new_n361), .A4(new_n491), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n588), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n301), .B2(new_n584), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n599), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n383), .A2(G264), .A3(G1698), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n383), .A2(G257), .A3(new_n281), .ZN(new_n609));
  INV_X1    g0409(.A(G303), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n280), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n289), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n458), .A2(G270), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n612), .A2(G190), .A3(new_n470), .A4(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n437), .B(new_n207), .C1(G33), .C2(new_n225), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G20), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n259), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n259), .A2(KEYINPUT20), .A3(new_n615), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n361), .A2(G116), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n492), .B2(G116), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n613), .A2(new_n470), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n301), .B1(new_n628), .B2(new_n612), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n607), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n612), .A2(new_n470), .A3(new_n613), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT87), .A3(new_n626), .A4(new_n614), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n307), .B1(new_n622), .B2(new_n624), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n628), .A2(new_n625), .A3(G179), .A4(new_n612), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n631), .B2(new_n638), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT88), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n634), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n606), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n434), .A2(new_n505), .A3(new_n576), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n316), .ZN(new_n650));
  INV_X1    g0450(.A(new_n336), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n374), .A2(new_n360), .B1(new_n379), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n432), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n427), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n654), .B2(new_n306), .ZN(new_n655));
  INV_X1    g0455(.A(new_n434), .ZN(new_n656));
  INV_X1    g0456(.A(new_n606), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n497), .A2(new_n498), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n473), .A2(new_n479), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n500), .B1(new_n660), .B2(KEYINPUT97), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n583), .A2(new_n289), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n301), .B1(new_n663), .B2(new_n579), .ZN(new_n664));
  INV_X1    g0464(.A(new_n603), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n589), .B(new_n665), .C1(new_n597), .C2(new_n265), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT94), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT94), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n604), .B(new_n668), .C1(new_n301), .C2(new_n584), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n669), .A3(new_n600), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n599), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n473), .A2(new_n479), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n661), .A2(new_n662), .A3(new_n672), .A4(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n659), .A2(new_n599), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n642), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n639), .A3(new_n640), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n557), .B1(new_n560), .B2(new_n312), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n555), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT96), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT96), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n643), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n671), .B1(new_n574), .B2(new_n570), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n499), .A2(new_n504), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(KEYINPUT95), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT95), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n499), .A2(new_n686), .A3(new_n689), .A4(new_n504), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n676), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n655), .B1(new_n656), .B2(new_n691), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n645), .A2(new_n647), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n693), .B1(new_n626), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n678), .A2(new_n625), .A3(new_n699), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n576), .B1(new_n567), .B2(new_n700), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n562), .B2(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n643), .A2(new_n699), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n576), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n680), .B2(new_n699), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT98), .ZN(G399));
  NOR2_X1   g0514(.A1(new_n210), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n594), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n217), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n648), .A2(new_n505), .A3(new_n576), .A4(new_n700), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n631), .A2(new_n312), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n450), .A2(new_n476), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n559), .A2(new_n514), .A3(new_n584), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n724), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n584), .B(KEYINPUT99), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n312), .A3(new_n560), .A4(new_n631), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n728), .B(new_n729), .C1(new_n503), .C2(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n699), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n722), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n687), .A2(KEYINPUT95), .ZN(new_n737));
  INV_X1    g0537(.A(new_n685), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n690), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n676), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n699), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n658), .A2(new_n662), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT100), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n501), .A2(new_n502), .A3(new_n471), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n724), .A2(G169), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT97), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n672), .A2(new_n747), .A3(new_n494), .A4(new_n674), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n744), .B1(new_n748), .B2(new_n662), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n747), .A2(new_n494), .A3(new_n674), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(KEYINPUT100), .A3(KEYINPUT26), .A4(new_n672), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n564), .A2(new_n565), .A3(new_n643), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n499), .A2(new_n753), .A3(new_n504), .A4(new_n686), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(new_n754), .A3(new_n599), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT29), .B(new_n700), .C1(new_n750), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n736), .B1(new_n742), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n720), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n209), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n206), .B1(new_n759), .B2(G45), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n716), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n705), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G330), .B2(new_n703), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n214), .B1(G20), .B2(new_n307), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n378), .A2(G179), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n207), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n225), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(KEYINPUT32), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n769), .B(new_n776), .C1(G87), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n207), .A2(new_n312), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n781), .A2(new_n301), .A3(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n781), .A2(new_n378), .A3(new_n301), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n231), .B1(new_n785), .B2(new_n202), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n780), .A2(new_n771), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(G77), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n770), .A2(new_n378), .A3(G200), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G107), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n781), .A2(new_n378), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G58), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n280), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(KEYINPUT32), .B2(new_n775), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n779), .A2(new_n789), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n318), .B1(new_n787), .B2(new_n799), .C1(new_n768), .C2(new_n512), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G303), .B2(new_n778), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n791), .A2(G283), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G326), .A2(new_n784), .B1(new_n782), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n772), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n793), .A2(G322), .B1(G329), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n766), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n765), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n406), .A2(new_n408), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n210), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n218), .A2(new_n462), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n462), .C2(new_n256), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n318), .A2(new_n210), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G355), .B1(new_n616), .B2(new_n210), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n808), .A2(new_n820), .A3(new_n761), .ZN(new_n821));
  INV_X1    g0621(.A(new_n811), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n703), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n764), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n651), .A2(new_n700), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n338), .B1(new_n333), .B2(new_n700), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n336), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n810), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n831), .A2(new_n783), .B1(new_n794), .B2(new_n512), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n785), .A2(new_n610), .B1(new_n772), .B2(new_n799), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n791), .A2(G87), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n778), .A2(G107), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n280), .B(new_n769), .C1(G116), .C2(new_n788), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n782), .A2(G150), .B1(G159), .B2(new_n788), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n785), .C1(new_n841), .C2(new_n794), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n791), .A2(G68), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n843), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n768), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G58), .B1(G132), .B2(new_n805), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(new_n814), .C1(new_n202), .C2(new_n777), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n838), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n765), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n765), .A2(new_n809), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(G77), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n762), .B1(new_n830), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT102), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n741), .B2(new_n829), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n741), .A2(new_n857), .A3(new_n829), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n339), .A2(new_n700), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n859), .A2(new_n860), .B1(new_n691), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(new_n736), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n761), .B1(new_n862), .B2(new_n736), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n856), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(KEYINPUT103), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  OR2_X1    g0669(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n215), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  NAND3_X1  g0673(.A1(new_n218), .A2(G77), .A3(new_n395), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n202), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n206), .B(G13), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n397), .B1(new_n411), .B2(new_n231), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n419), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n259), .A3(new_n412), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n394), .B1(new_n881), .B2(new_n425), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n421), .A2(new_n425), .A3(new_n430), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT104), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n412), .A2(new_n259), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n424), .B1(new_n886), .B2(new_n880), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n431), .C1(new_n887), .C2(new_n394), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n697), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n421), .A2(new_n425), .ZN(new_n891));
  INV_X1    g0691(.A(new_n697), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT105), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT105), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n894), .B(new_n697), .C1(new_n421), .C2(new_n425), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n883), .A2(new_n426), .A3(KEYINPUT37), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n890), .A2(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n889), .B1(new_n427), .B2(new_n432), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n883), .A2(new_n426), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n893), .B2(new_n895), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n893), .A2(new_n895), .ZN(new_n906));
  INV_X1    g0706(.A(new_n426), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n431), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n905), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n897), .B(KEYINPUT106), .C1(new_n893), .C2(new_n895), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n433), .A2(new_n906), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n878), .B1(new_n901), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n916));
  INV_X1    g0716(.A(new_n900), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n887), .A2(new_n697), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n431), .B1(new_n887), .B2(new_n394), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(KEYINPUT104), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n908), .B1(new_n920), .B2(new_n888), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n902), .B(new_n908), .C1(new_n893), .C2(new_n895), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT38), .B(new_n917), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n916), .A2(new_n924), .A3(KEYINPUT39), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n375), .A2(new_n699), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n374), .A2(new_n699), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n375), .A2(new_n379), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n375), .B2(new_n379), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n861), .B1(new_n739), .B2(new_n740), .ZN(new_n934));
  INV_X1    g0734(.A(new_n826), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n916), .A2(new_n924), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n427), .A2(new_n892), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n928), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n434), .B(new_n756), .C1(new_n741), .C2(KEYINPUT29), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n655), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n940), .B(new_n942), .Z(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n829), .B1(new_n930), .B2(new_n931), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n722), .B2(new_n735), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n946), .B2(KEYINPUT107), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT108), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n901), .B2(new_n914), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n896), .B1(new_n427), .B2(new_n432), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n922), .A2(new_n905), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n911), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n924), .B(KEYINPUT108), .C1(new_n954), .C2(KEYINPUT38), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n947), .A2(new_n949), .A3(new_n951), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n946), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n948), .B1(new_n957), .B2(new_n937), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n722), .A2(new_n735), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n434), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n959), .A2(new_n961), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n962), .A2(new_n963), .A3(new_n721), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n944), .A2(new_n964), .B1(new_n206), .B2(new_n759), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n944), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n877), .B1(new_n965), .B2(new_n966), .ZN(G367));
  OAI211_X1 g0767(.A(new_n499), .B(new_n504), .C1(new_n500), .C2(new_n700), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n751), .A2(new_n699), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n968), .A2(KEYINPUT111), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT111), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n708), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n666), .A2(new_n699), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n672), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n599), .B2(new_n974), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(KEYINPUT109), .B2(new_n975), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT110), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n972), .A2(new_n711), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT42), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n566), .B1(new_n970), .B2(new_n971), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n699), .B1(new_n983), .B2(new_n499), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(KEYINPUT43), .A2(new_n980), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n988), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n973), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT112), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n973), .A3(new_n990), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n715), .B(KEYINPUT41), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n972), .A2(new_n712), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT44), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n972), .A2(new_n712), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT45), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n997), .A2(new_n708), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n708), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n711), .B1(new_n707), .B2(new_n710), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(new_n704), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n757), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n995), .B1(new_n1006), .B2(new_n757), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n760), .B(KEYINPUT113), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n994), .B1(new_n992), .B2(new_n993), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n815), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n812), .B1(new_n211), .B2(new_n327), .C1(new_n1011), .C2(new_n247), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1012), .A2(new_n762), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n848), .A2(G68), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n794), .B2(new_n268), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n805), .A2(G137), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n782), .A2(G159), .B1(new_n784), .B2(G143), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n280), .B1(new_n787), .B2(new_n202), .C1(new_n795), .C2(new_n777), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n790), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(G77), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n794), .A2(new_n610), .B1(new_n785), .B2(new_n799), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G97), .B2(new_n1020), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n814), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n480), .C2(new_n768), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n782), .A2(G294), .B1(G283), .B2(new_n788), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n777), .B2(new_n616), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n805), .A2(G317), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1022), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n1013), .B1(new_n766), .B2(new_n1034), .C1(new_n980), .C2(new_n822), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1010), .A2(new_n1035), .ZN(G387));
  NOR2_X1   g0836(.A1(new_n1005), .A2(new_n757), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1005), .A2(new_n757), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n715), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n818), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1041), .A2(new_n717), .B1(G107), .B2(new_n211), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n244), .A2(new_n462), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n717), .B(new_n462), .C1(new_n231), .C2(new_n283), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n266), .B2(G50), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n324), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1011), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n762), .B1(new_n1050), .B2(new_n813), .ZN(new_n1051));
  INV_X1    g0851(.A(G326), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n790), .A2(new_n616), .B1(new_n772), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n793), .A2(G317), .B1(new_n784), .B2(G322), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n782), .A2(G311), .B1(G303), .B2(new_n788), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n768), .A2(new_n831), .B1(new_n777), .B2(new_n512), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n814), .B(new_n1053), .C1(new_n1060), .C2(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT49), .B2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n783), .A2(new_n266), .B1(new_n785), .B2(new_n773), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n794), .A2(new_n202), .B1(new_n787), .B2(new_n231), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n768), .A2(new_n327), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n777), .A2(new_n283), .B1(new_n772), .B2(new_n268), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT115), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n791), .A2(G97), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n814), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1051), .B1(new_n1072), .B2(new_n765), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n707), .B2(new_n822), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1040), .A2(new_n1076), .ZN(G393));
  OAI21_X1  g0877(.A(new_n1039), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1006), .A2(new_n715), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n793), .A2(G311), .B1(new_n784), .B2(G317), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  OAI21_X1  g0881(.A(new_n318), .B1(new_n787), .B2(new_n512), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n783), .A2(new_n610), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G322), .C2(new_n805), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n848), .A2(G116), .B1(new_n778), .B2(G283), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1084), .A3(new_n792), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n787), .A2(new_n266), .B1(new_n772), .B2(new_n841), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G50), .B2(new_n782), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n768), .A2(new_n283), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G68), .B2(new_n778), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1090), .A3(new_n814), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n793), .A2(G159), .B1(new_n784), .B2(G150), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n835), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n765), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n253), .A2(new_n815), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n812), .B1(new_n225), .B2(new_n211), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n762), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n972), .B2(new_n811), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1079), .A2(new_n1101), .ZN(G390));
  AND3_X1   g0902(.A1(new_n736), .A2(new_n829), .A3(new_n933), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n927), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n951), .A2(new_n1104), .A3(new_n955), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n700), .B(new_n828), .C1(new_n750), .C2(new_n755), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n932), .B1(new_n1106), .B2(new_n826), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n936), .A2(new_n1104), .B1(new_n915), .B2(new_n925), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n736), .A2(new_n829), .A3(new_n933), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n826), .B1(new_n691), .B2(new_n861), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n927), .B1(new_n1112), .B2(new_n933), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1111), .B1(new_n1105), .B2(new_n1107), .C1(new_n926), .C2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1114), .A3(new_n1009), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT118), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n761), .B1(new_n266), .B2(new_n853), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n783), .A2(new_n840), .B1(new_n787), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G159), .B2(new_n848), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n778), .A2(G150), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n793), .A2(G132), .B1(G125), .B2(new_n805), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n280), .C1(new_n1126), .C2(new_n785), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1124), .B(new_n1127), .C1(G50), .C2(new_n1020), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n783), .A2(new_n480), .B1(new_n785), .B2(new_n831), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n794), .A2(new_n616), .B1(new_n787), .B2(new_n225), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n318), .B1(new_n772), .B2(new_n512), .C1(new_n223), .C2(new_n777), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1089), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1122), .A2(new_n1128), .B1(new_n845), .B2(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1118), .B1(new_n766), .B2(new_n1133), .C1(new_n926), .C2(new_n810), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1117), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n434), .A2(new_n736), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n941), .A2(new_n655), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n933), .B1(new_n736), .B2(new_n829), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1112), .B1(new_n1103), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n960), .A2(G330), .A3(new_n829), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n932), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(new_n826), .A3(new_n1111), .A4(new_n1106), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1110), .A2(new_n1114), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT116), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1110), .A2(new_n1114), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(KEYINPUT117), .A3(new_n715), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n716), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT117), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1136), .B1(new_n1153), .B2(new_n1155), .ZN(G378));
  NAND3_X1  g0956(.A1(new_n956), .A2(G330), .A3(new_n958), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n306), .A2(new_n316), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n273), .A2(new_n892), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT122), .Z(new_n1162));
  XNOR2_X1  g0962(.A(new_n1160), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n956), .A2(G330), .A3(new_n958), .A4(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n940), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n940), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(new_n809), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n848), .A2(G150), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n777), .A2(new_n1119), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT120), .Z(new_n1175));
  AOI22_X1  g0975(.A1(new_n782), .A2(G132), .B1(new_n784), .B2(G125), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n793), .A2(G128), .B1(G137), .B2(new_n788), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1020), .A2(G159), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1184), .B2(new_n1178), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1014), .B1(new_n783), .B2(new_n225), .C1(new_n480), .C2(new_n794), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1025), .A2(new_n452), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n587), .A2(new_n788), .B1(new_n805), .B2(G283), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n616), .B2(new_n785), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n795), .A2(new_n790), .B1(new_n777), .B2(new_n283), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1187), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n765), .B1(new_n1185), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT121), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n761), .B(new_n1197), .C1(new_n202), .C2(new_n853), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1171), .A2(new_n1009), .B1(new_n1172), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1138), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n715), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1138), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1149), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1171), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1199), .B1(new_n1204), .B2(new_n1207), .ZN(G375));
  NAND2_X1  g1008(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1205), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1140), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n995), .B(KEYINPUT123), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n932), .A2(new_n809), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n762), .B1(G68), .B2(new_n854), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n616), .A2(new_n783), .B1(new_n794), .B2(new_n831), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n785), .A2(new_n512), .B1(new_n772), .B2(new_n610), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n791), .A2(G77), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n778), .A2(G97), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n280), .B(new_n1065), .C1(G107), .C2(new_n788), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n784), .A2(G132), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n794), .B2(new_n840), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G58), .B2(new_n1020), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n783), .A2(new_n1119), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G150), .A2(new_n788), .B1(new_n805), .B2(G128), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n848), .A2(G50), .B1(new_n778), .B2(G159), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1229), .B2(new_n1025), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n766), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1215), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1209), .A2(new_n1009), .B1(new_n1214), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1213), .A2(new_n1235), .ZN(G381));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1079), .A2(new_n1101), .A3(new_n1237), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G387), .A2(G384), .A3(G381), .A4(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1154), .A2(KEYINPUT117), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1151), .B1(new_n1154), .B2(KEYINPUT117), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1135), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1172), .A2(new_n1198), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1008), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n716), .B1(new_n1206), .B2(new_n1201), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1200), .B1(new_n1244), .B2(new_n1203), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1239), .A2(new_n1242), .A3(new_n1248), .ZN(G407));
  NAND2_X1  g1049(.A1(new_n698), .A2(G213), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(new_n1242), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  XNOR2_X1  g1053(.A(G393), .B(new_n824), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(G390), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(G390), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1010), .A2(new_n1255), .A3(new_n1035), .A4(new_n1256), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1248), .A2(G378), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1206), .A2(new_n1171), .A3(new_n1212), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1199), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1242), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1251), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1210), .A2(KEYINPUT60), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1211), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n716), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1267), .B2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1235), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n868), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT62), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1250), .ZN(new_n1276));
  AOI211_X1 g1076(.A(KEYINPUT125), .B(new_n1251), .C1(new_n1261), .C2(new_n1264), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1273), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1251), .A2(G2897), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1271), .B(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1260), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1272), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1265), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1271), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1260), .A2(KEYINPUT61), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1287), .A2(new_n1290), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1293), .ZN(G405));
  NOR2_X1   g1094(.A1(G375), .A2(new_n1242), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1248), .A2(G378), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1271), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1242), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1272), .A2(new_n1298), .A3(new_n1261), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT127), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1260), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1297), .A2(new_n1299), .A3(KEYINPUT126), .A4(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1302), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1302), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(G402));
endmodule


