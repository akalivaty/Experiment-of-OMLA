//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n212), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n210), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G58), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XNOR2_X1  g0041(.A(KEYINPUT3), .B(G33), .ZN(new_n242));
  AND2_X1   g0042(.A1(new_n242), .A2(G1698), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n243), .A2(G223), .B1(G77), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G222), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n251), .A2(new_n245), .A3(new_n247), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n258), .B(G274), .C1(G41), .C2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(G226), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G200), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n246), .A2(G20), .ZN(new_n268));
  XOR2_X1   g0068(.A(KEYINPUT8), .B(G58), .Z(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  INV_X1    g0070(.A(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n246), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n268), .A2(new_n269), .B1(new_n274), .B2(G150), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n271), .B2(new_n202), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n255), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(new_n258), .B2(G20), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G50), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n266), .A2(new_n267), .B1(new_n285), .B2(KEYINPUT9), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n257), .A2(new_n265), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n288), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(new_n291), .B(KEYINPUT10), .Z(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n285), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n266), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n295), .B2(new_n294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n245), .A2(new_n247), .A3(G232), .A4(G1698), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n302), .C1(new_n253), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n256), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n262), .A2(G238), .A3(new_n263), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n259), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT13), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n288), .ZN(new_n314));
  INV_X1    g0114(.A(new_n274), .ZN(new_n315));
  INV_X1    g0115(.A(G50), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n268), .A2(G77), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n271), .B2(G68), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n278), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT11), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n280), .A2(KEYINPUT12), .A3(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT12), .B1(new_n280), .B2(G68), .ZN(new_n325));
  AOI22_X1  g0125(.A1(G68), .A2(new_n282), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n314), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n313), .A2(KEYINPUT71), .A3(G200), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT71), .B1(new_n313), .B2(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n311), .B1(new_n305), .B2(new_n308), .ZN(new_n333));
  AOI211_X1 g0133(.A(KEYINPUT13), .B(new_n307), .C1(new_n304), .C2(new_n256), .ZN(new_n334));
  OAI21_X1  g0134(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT14), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(G169), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n310), .A2(G179), .A3(new_n312), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n327), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n251), .A2(G223), .A3(new_n252), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G226), .A2(G1698), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n248), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n246), .A2(new_n217), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n256), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT74), .A4(G232), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n260), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n352), .A3(new_n288), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n347), .A2(new_n352), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G200), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT73), .B1(new_n244), .B2(G33), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n246), .A3(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n359), .A3(new_n245), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n242), .B2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n212), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G58), .A2(G68), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G58), .A3(G68), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(new_n213), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n274), .A2(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n356), .B1(new_n365), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n248), .B2(new_n271), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n361), .B(G20), .C1(new_n245), .C2(new_n247), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(G20), .A2(new_n370), .B1(new_n274), .B2(G159), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n278), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n269), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n258), .B2(G20), .ZN(new_n382));
  INV_X1    g0182(.A(new_n280), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n278), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n382), .A2(new_n384), .B1(new_n383), .B2(new_n381), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n355), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n385), .ZN(new_n389));
  INV_X1    g0189(.A(new_n278), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n271), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n212), .B1(new_n364), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n373), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n389), .B1(new_n394), .B2(new_n374), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT17), .B1(new_n395), .B2(new_n355), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n380), .A2(new_n385), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n347), .A2(new_n352), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G169), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n347), .A2(new_n352), .A3(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT18), .B1(new_n399), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT15), .B(G87), .Z(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n315), .B2(new_n381), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n278), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n280), .A2(G77), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n282), .B2(G77), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n264), .A2(G244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n259), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n243), .A2(G238), .B1(G107), .B2(new_n248), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT66), .B(G1698), .Z(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n242), .A3(G232), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n420), .B2(new_n256), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n414), .B1(new_n422), .B2(new_n293), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n421), .A2(KEYINPUT70), .A3(new_n296), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT70), .B1(new_n421), .B2(new_n296), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n421), .B2(new_n267), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n414), .B(KEYINPUT69), .C1(new_n267), .C2(new_n421), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(G190), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n427), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n300), .A2(new_n342), .A3(new_n407), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n244), .A2(G33), .ZN(new_n438));
  OAI21_X1  g0238(.A(G303), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n245), .A2(new_n247), .A3(G264), .A4(G1698), .ZN(new_n440));
  INV_X1    g0240(.A(G257), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n439), .B(new_n440), .C1(new_n253), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n418), .A2(new_n242), .A3(G257), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT80), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n440), .A4(new_n439), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n446), .A3(new_n256), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n262), .A2(G274), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n256), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(G270), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n447), .A2(KEYINPUT81), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT81), .B1(new_n447), .B2(new_n457), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n458), .A2(new_n459), .A3(new_n267), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n280), .A2(G116), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n384), .B1(G1), .B2(new_n246), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n271), .C1(G33), .C2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n278), .C1(new_n271), .C2(G116), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n436), .B1(new_n460), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n447), .A2(new_n457), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n447), .A2(KEYINPUT81), .A3(new_n457), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT82), .B(new_n471), .C1(new_n478), .C2(new_n267), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(G190), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n262), .B(G250), .C1(G1), .C2(new_n449), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n450), .A2(G274), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n242), .A2(G244), .A3(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n216), .C2(new_n253), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n487), .B2(new_n256), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n293), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n296), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n245), .A2(new_n247), .A3(new_n271), .A4(G68), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT77), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n242), .A2(KEYINPUT77), .A3(new_n271), .A4(G68), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n271), .A2(G33), .A3(G97), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n271), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT76), .ZN(new_n503));
  INV_X1    g0303(.A(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n217), .A2(new_n466), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n502), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n278), .B1(new_n500), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n408), .A2(new_n280), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n463), .A2(new_n408), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n492), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n489), .A2(new_n288), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n489), .A2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n463), .A2(G87), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n493), .A2(new_n494), .B1(new_n498), .B2(new_n497), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(new_n496), .C1(new_n506), .C2(new_n507), .ZN(new_n523));
  AOI211_X1 g0323(.A(KEYINPUT78), .B(new_n510), .C1(new_n523), .C2(new_n278), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n514), .B1(new_n509), .B2(new_n511), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n520), .B(new_n521), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n516), .A2(KEYINPUT79), .A3(new_n520), .A4(new_n521), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n518), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n293), .B1(new_n464), .B2(new_n470), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n476), .A2(new_n477), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n476), .A2(KEYINPUT21), .A3(new_n477), .A4(new_n531), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n447), .A2(G179), .A3(new_n457), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n471), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n245), .A2(new_n247), .A3(G257), .A4(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n253), .C2(new_n218), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n256), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n455), .A2(G274), .A3(new_n262), .A4(new_n450), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n456), .A2(G264), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n293), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n543), .A2(new_n256), .B1(G264), .B2(new_n456), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n296), .A3(new_n545), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n383), .A2(KEYINPUT25), .A3(new_n504), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n280), .B2(G107), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n462), .B2(new_n504), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n245), .A2(new_n247), .A3(new_n271), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT22), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n242), .A2(new_n559), .A3(new_n271), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n271), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n504), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n271), .A2(G33), .A3(G116), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n390), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n558), .B2(new_n560), .ZN(new_n574));
  INV_X1    g0374(.A(new_n572), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n556), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n540), .B1(new_n551), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n544), .A2(new_n288), .A3(new_n545), .A4(new_n546), .ZN(new_n579));
  AOI221_X4 g0379(.A(new_n454), .B1(new_n456), .B2(G264), .C1(new_n543), .C2(new_n256), .ZN(new_n580));
  OAI211_X1 g0380(.A(KEYINPUT85), .B(new_n579), .C1(new_n580), .C2(G200), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n579), .A2(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n556), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n278), .B1(new_n574), .B2(new_n575), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n571), .A2(new_n572), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(KEYINPUT84), .A3(new_n550), .A4(new_n548), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n578), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n590), .A2(new_n466), .A3(G107), .ZN(new_n591));
  XNOR2_X1  g0391(.A(G97), .B(G107), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n593), .A2(new_n271), .B1(new_n203), .B2(new_n315), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n504), .B1(new_n363), .B2(new_n364), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n278), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n280), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n463), .B2(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n453), .A2(new_n262), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n545), .B1(new_n601), .B2(new_n441), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  INV_X1    g0403(.A(G244), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n253), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n418), .A2(new_n242), .A3(KEYINPUT4), .A4(G244), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n242), .A2(G250), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n465), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n602), .B1(new_n608), .B2(new_n256), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G190), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT75), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI211_X1 g0412(.A(KEYINPUT75), .B(new_n602), .C1(new_n608), .C2(new_n256), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n600), .B(new_n610), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n609), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n293), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n296), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n599), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n589), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n481), .A2(new_n530), .A3(new_n539), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n435), .A2(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n332), .A2(new_n427), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n398), .B1(new_n623), .B2(new_n341), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n404), .B2(new_n405), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT18), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n293), .B1(new_n347), .B2(new_n352), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G179), .B2(new_n354), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n395), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(KEYINPUT88), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n292), .B1(new_n624), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n298), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT86), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(KEYINPUT86), .B(new_n521), .C1(new_n524), .C2(new_n525), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n519), .B1(G200), .B2(new_n489), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n518), .ZN(new_n643));
  INV_X1    g0443(.A(new_n618), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n530), .A2(new_n644), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n551), .A2(new_n577), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n537), .B1(new_n532), .B2(new_n533), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT87), .A3(new_n535), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n614), .A2(new_n583), .A3(new_n618), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n643), .A3(new_n641), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n646), .B(new_n648), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n635), .B1(new_n435), .B2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n458), .A2(new_n459), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n288), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n472), .B1(new_n662), .B2(G200), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(KEYINPUT82), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n650), .B1(new_n665), .B2(new_n473), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n258), .A2(new_n271), .A3(G13), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n670));
  INV_X1    g0470(.A(G213), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(G343), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT90), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n666), .B1(new_n471), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n652), .A2(new_n472), .A3(new_n654), .A4(new_n679), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n661), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n589), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n577), .B2(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n649), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n539), .A2(new_n679), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n689), .A2(new_n684), .B1(new_n649), .B2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(G399));
  NOR2_X1   g0491(.A1(new_n505), .A2(G116), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G41), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n207), .A2(KEYINPUT92), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT92), .B1(new_n207), .B2(new_n695), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n694), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n214), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n666), .A2(new_n530), .A3(new_n620), .A4(new_n680), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n580), .A2(G179), .A3(new_n488), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n476), .A3(new_n477), .A4(new_n615), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n488), .A2(new_n549), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n609), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n536), .ZN(new_n710));
  INV_X1    g0510(.A(new_n536), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n609), .A4(new_n708), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n679), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(new_n679), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n661), .B1(new_n704), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n653), .A2(new_n535), .A3(new_n578), .A4(new_n588), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n643), .A3(new_n641), .A4(new_n656), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n528), .A2(new_n529), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n723), .A3(new_n643), .A4(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT93), .A3(new_n680), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT93), .B1(new_n726), .B2(new_n680), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n658), .A2(new_n680), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n719), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n703), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n258), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n699), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n683), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n681), .A2(new_n682), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(G330), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n255), .B1(G20), .B2(new_n293), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n271), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n296), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n267), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n748), .A2(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n271), .A2(new_n288), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n242), .B(new_n753), .C1(G303), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n296), .A2(new_n267), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n745), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n760), .A2(G326), .B1(new_n763), .B2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(new_n754), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(new_n296), .A3(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n758), .A2(new_n745), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G322), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G294), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n757), .A2(new_n764), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n748), .A2(KEYINPUT96), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G77), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n242), .B1(new_n780), .B2(new_n211), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G97), .B2(new_n772), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n762), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n759), .A2(new_n316), .B1(new_n755), .B2(new_n217), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n767), .A2(new_n212), .B1(new_n751), .B2(new_n504), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n779), .A2(new_n782), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n744), .B1(new_n774), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n743), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  NAND2_X1  g0595(.A1(new_n237), .A2(G45), .ZN(new_n796));
  INV_X1    g0596(.A(new_n207), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n242), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G45), .C2(new_n214), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n242), .A2(new_n207), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(G116), .B2(new_n207), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  AOI21_X1  g0603(.A(new_n795), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n739), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n790), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n793), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n741), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n742), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  OAI211_X1 g0610(.A(new_n423), .B(new_n680), .C1(new_n425), .C2(new_n424), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n680), .A2(new_n414), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n433), .B2(new_n430), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n813), .B2(new_n427), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n730), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n811), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n433), .A2(new_n430), .ZN(new_n817));
  INV_X1    g0617(.A(new_n812), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(new_n819), .B2(new_n426), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n658), .A2(new_n680), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n718), .B1(new_n621), .B2(new_n679), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G330), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n739), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n824), .B2(new_n822), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n743), .A2(new_n791), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n805), .B1(new_n203), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G107), .A2(new_n756), .B1(new_n768), .B2(G283), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n749), .B2(new_n762), .ZN(new_n830));
  INV_X1    g0630(.A(new_n751), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n766), .A2(G294), .B1(G87), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n242), .B1(new_n760), .B2(G303), .ZN(new_n833));
  INV_X1    g0633(.A(new_n772), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n833), .C1(new_n466), .C2(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n830), .B(new_n835), .C1(new_n778), .C2(G116), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n211), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G50), .A2(new_n756), .B1(new_n763), .B2(G132), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n242), .C1(new_n212), .C2(new_n751), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n766), .A2(G143), .B1(new_n760), .B2(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n767), .C1(new_n777), .C2(new_n783), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n837), .B(new_n839), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n836), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n828), .B1(new_n744), .B2(new_n846), .C1(new_n820), .C2(new_n792), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n826), .A2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(G116), .ZN(new_n849));
  INV_X1    g0649(.A(new_n593), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n849), .B(new_n210), .C1(new_n850), .C2(KEYINPUT35), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(KEYINPUT35), .B2(new_n850), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n367), .A2(new_n369), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n213), .A2(G50), .A3(G77), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(G50), .B2(new_n212), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(G1), .A3(new_n735), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT97), .Z(new_n859));
  NAND3_X1  g0659(.A1(new_n626), .A2(new_n397), .A3(new_n632), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n399), .A2(new_n674), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n625), .B1(new_n395), .B2(new_n629), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  AOI21_X1  g0665(.A(G200), .B1(new_n347), .B2(new_n352), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n288), .B2(new_n354), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n399), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n861), .B1(new_n386), .B2(new_n865), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n399), .B2(new_n867), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n629), .A2(new_n673), .B1(new_n380), .B2(new_n385), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT99), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n401), .A2(new_n402), .A3(new_n673), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n399), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT99), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n386), .A4(new_n873), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n356), .B1(new_n392), .B2(new_n373), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n379), .A2(new_n886), .A3(new_n278), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n385), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n674), .B(new_n888), .C1(new_n398), .C2(new_n406), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n877), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n873), .B1(new_n891), .B2(new_n386), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n881), .B2(new_n893), .ZN(new_n894));
  AOI211_X1 g0694(.A(KEYINPUT100), .B(new_n892), .C1(new_n876), .C2(new_n880), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n889), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n885), .A2(new_n896), .A3(KEYINPUT102), .ZN(new_n897));
  INV_X1    g0697(.A(new_n880), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n395), .B2(new_n355), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n879), .B1(new_n899), .B2(new_n878), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n893), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT100), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n881), .A2(new_n890), .A3(new_n893), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT38), .A4(new_n889), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n337), .B1(new_n313), .B2(G169), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n338), .A2(new_n339), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n327), .B(new_n679), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT98), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT98), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n340), .A2(new_n912), .A3(new_n327), .A4(new_n679), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n679), .A2(new_n327), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n332), .A2(new_n341), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n820), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n704), .B2(new_n718), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n884), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n896), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n919), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n907), .A2(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n435), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n925), .A2(new_n926), .A3(new_n823), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n823), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n927), .A2(new_n928), .A3(new_n661), .ZN(new_n929));
  INV_X1    g0729(.A(new_n917), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n821), .B2(new_n811), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n922), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n897), .A2(new_n933), .A3(new_n906), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n340), .A2(new_n327), .A3(new_n680), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n921), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n633), .A2(new_n673), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n729), .A2(new_n926), .A3(new_n732), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n635), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n929), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n258), .B2(new_n736), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n929), .A2(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n859), .B1(new_n945), .B2(new_n946), .ZN(G367));
  INV_X1    g0747(.A(new_n733), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  INV_X1    g0750(.A(new_n619), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n679), .A2(new_n599), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(new_n952), .B1(new_n644), .B2(new_n679), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n690), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n950), .B1(new_n690), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n689), .A2(new_n684), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n649), .A2(new_n680), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT105), .B1(new_n960), .B2(new_n953), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n690), .A2(new_n950), .A3(new_n954), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(KEYINPUT44), .A3(new_n953), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n690), .B2(new_n954), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n688), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n957), .A2(new_n963), .A3(new_n688), .A4(new_n967), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n958), .B1(new_n687), .B2(new_n689), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n741), .A2(G330), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT107), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT106), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT107), .B1(new_n683), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(KEYINPUT107), .B(new_n973), .C1(new_n683), .C2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n948), .B1(new_n972), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n699), .B(KEYINPUT41), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n737), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n954), .A2(new_n684), .A3(new_n689), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n985), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT104), .B1(new_n985), .B2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n578), .A2(new_n588), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n614), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n679), .B1(new_n989), .B2(new_n618), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n985), .B2(KEYINPUT42), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n680), .B1(new_n638), .B2(new_n639), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n518), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n641), .A2(new_n643), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n993), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT103), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(KEYINPUT103), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n992), .B(new_n1001), .C1(new_n999), .C2(new_n997), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n992), .B2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n688), .A2(new_n953), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n984), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n408), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n798), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n794), .B1(new_n207), .B2(new_n1007), .C1(new_n232), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n739), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT108), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n242), .B1(new_n751), .B2(new_n203), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n777), .A2(new_n316), .B1(KEYINPUT109), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(KEYINPUT109), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n772), .A2(G68), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n211), .B2(new_n755), .C1(new_n780), .C2(new_n841), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G143), .A2(new_n760), .B1(new_n768), .B2(G159), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n762), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n751), .A2(new_n466), .B1(new_n762), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(G303), .ZN(new_n1023));
  INV_X1    g0823(.A(G294), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n780), .A2(new_n1023), .B1(new_n767), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(new_n778), .C2(G283), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n248), .B1(new_n759), .B2(new_n749), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n756), .A2(G116), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(new_n834), .B2(new_n504), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1027), .B(new_n1030), .C1(new_n1029), .C2(new_n1028), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1014), .A2(new_n1020), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT110), .Z(new_n1033));
  INV_X1    g0833(.A(KEYINPUT47), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n743), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1011), .B1(new_n807), .B2(new_n996), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1006), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(G387));
  NAND3_X1  g0840(.A1(new_n685), .A2(new_n686), .A3(new_n793), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n798), .B1(new_n229), .B2(new_n449), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n694), .B2(new_n800), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n269), .A2(new_n316), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT50), .Z(new_n1045));
  AOI21_X1  g0845(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n694), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1043), .A2(new_n1047), .B1(new_n504), .B2(new_n797), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n739), .B1(new_n1048), .B2(new_n795), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n747), .A2(G68), .B1(new_n768), .B2(new_n269), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n834), .A2(new_n1007), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n248), .B(new_n1052), .C1(G97), .C2(new_n831), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n755), .A2(new_n203), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G159), .B2(new_n760), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n766), .A2(G50), .B1(G150), .B2(new_n763), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n242), .B1(new_n763), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n834), .A2(new_n752), .B1(new_n755), .B2(new_n1024), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G322), .A2(new_n760), .B1(new_n768), .B2(G311), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1021), .B2(new_n780), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n778), .B2(G303), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1058), .B1(new_n849), .B2(new_n751), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1049), .B1(new_n1068), .B2(new_n743), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n981), .A2(new_n738), .B1(new_n1041), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n981), .A2(new_n733), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n699), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n981), .A2(new_n733), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1071), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n700), .B1(new_n1075), .B2(new_n972), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT113), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n970), .A2(new_n971), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n1071), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1079), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n699), .B1(new_n1078), .B2(new_n1071), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT113), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n240), .A2(new_n798), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n794), .B1(new_n466), .B2(new_n207), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n766), .A2(G159), .B1(new_n760), .B2(G150), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n763), .A2(G143), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n316), .B2(new_n767), .C1(new_n212), .C2(new_n755), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n772), .A2(G77), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n242), .C1(new_n217), .C2(new_n751), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n778), .C2(new_n269), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n248), .B1(new_n751), .B2(new_n504), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G283), .A2(new_n756), .B1(new_n763), .B2(G322), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n1023), .B2(new_n767), .C1(new_n1024), .C2(new_n748), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G116), .C2(new_n772), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n766), .A2(G311), .B1(new_n760), .B2(G317), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n1087), .A2(new_n1092), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n739), .B1(new_n1084), .B2(new_n1085), .C1(new_n1099), .C2(new_n744), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n953), .B2(new_n793), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1078), .A2(KEYINPUT112), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n737), .B1(new_n1078), .B2(KEYINPUT112), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1080), .A2(new_n1083), .A3(new_n1104), .ZN(G390));
  NOR2_X1   g0905(.A1(new_n824), .A2(new_n918), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n897), .A2(new_n935), .A3(new_n906), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n819), .A2(new_n426), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n727), .B2(new_n728), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n811), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1110), .B2(new_n917), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n821), .A2(new_n811), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n917), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1113), .A2(new_n935), .B1(new_n937), .B2(new_n934), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1106), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n934), .A2(new_n937), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n931), .B2(new_n936), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n814), .B1(new_n916), .B2(new_n914), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n719), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n930), .B1(new_n1109), .B2(new_n811), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1119), .C1(new_n1120), .C2(new_n1107), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1115), .A2(new_n738), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n791), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n805), .B1(new_n381), .B2(new_n827), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n778), .A2(G97), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n751), .A2(new_n212), .B1(new_n762), .B2(new_n1024), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n242), .B(new_n1126), .C1(G87), .C2(new_n756), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n780), .A2(new_n849), .B1(new_n767), .B2(new_n504), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G283), .B2(new_n760), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1125), .A2(new_n1090), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n766), .A2(G132), .B1(G125), .B2(new_n763), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G128), .A2(new_n760), .B1(new_n768), .B2(G137), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n783), .C2(new_n834), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n242), .B1(new_n751), .B2(new_n316), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT116), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n755), .A2(new_n841), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1135), .B(new_n1137), .C1(new_n777), .C2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1130), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(KEYINPUT117), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(KEYINPUT117), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n743), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1123), .B(new_n1124), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1122), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1122), .A2(KEYINPUT118), .A3(new_n1144), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n930), .B1(new_n824), .B2(new_n814), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1151), .A2(new_n1119), .B1(new_n811), .B2(new_n821), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n726), .A2(new_n680), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT93), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n726), .A2(KEYINPUT93), .A3(new_n680), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n816), .B1(new_n1157), .B2(new_n1108), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n917), .B1(new_n719), .B2(new_n820), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n1106), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1152), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n926), .A2(new_n719), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n941), .A2(new_n635), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT114), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT114), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1109), .A2(new_n811), .A3(new_n1119), .A4(new_n1151), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1112), .B1(new_n1159), .B2(new_n1106), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1150), .A2(new_n1164), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1115), .A2(new_n1172), .A3(new_n1121), .ZN(new_n1173));
  AND4_X1   g0973(.A1(KEYINPUT115), .A2(new_n1171), .A3(new_n699), .A4(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1173), .A2(new_n699), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT115), .B1(new_n1175), .B2(new_n1171), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1149), .B1(new_n1174), .B2(new_n1176), .ZN(G378));
  NAND4_X1  g0977(.A1(new_n897), .A2(new_n919), .A3(KEYINPUT40), .A4(new_n906), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n823), .A2(new_n1118), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n921), .B2(new_n896), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(G330), .C1(KEYINPUT40), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT121), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n923), .A2(new_n924), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1184), .A2(KEYINPUT121), .A3(G330), .A4(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n284), .A2(new_n674), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n299), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1188), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1187), .B(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n925), .A2(new_n1192), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n940), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n940), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1190), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n738), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n805), .B1(new_n316), .B2(new_n827), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n747), .A2(new_n408), .B1(new_n768), .B2(G97), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT119), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G58), .A2(new_n831), .B1(new_n763), .B2(G283), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n849), .B2(new_n759), .C1(new_n504), .C2(new_n780), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1054), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n695), .A3(new_n248), .A4(new_n1015), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT120), .Z(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n748), .A2(new_n1018), .B1(new_n755), .B2(new_n1138), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G125), .A2(new_n760), .B1(new_n768), .B2(G132), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n841), .B2(new_n834), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G128), .C2(new_n766), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n783), .B2(new_n751), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n695), .B1(new_n244), .B2(new_n246), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1216), .A2(new_n1219), .B1(new_n316), .B2(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1209), .A2(new_n1210), .A3(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1199), .B1(new_n744), .B2(new_n1222), .C1(new_n1189), .C2(new_n792), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1198), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1173), .A2(new_n1165), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n699), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1190), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1196), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1173), .A2(new_n1165), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1227), .B2(new_n1232), .ZN(G375));
  INV_X1    g1033(.A(new_n983), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1170), .A2(new_n1164), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT122), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n805), .B1(new_n212), .B2(new_n827), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n766), .A2(G283), .B1(G97), .B2(new_n756), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1024), .B2(new_n759), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n778), .B2(G107), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n248), .B1(new_n751), .B2(new_n203), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n767), .A2(new_n849), .B1(new_n762), .B2(new_n1023), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1052), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n242), .B1(new_n751), .B2(new_n211), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n760), .A2(G132), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n780), .B2(new_n1018), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(G50), .C2(new_n772), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n767), .A2(new_n1138), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n748), .A2(new_n841), .B1(new_n783), .B2(new_n755), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G128), .C2(new_n763), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1241), .A2(new_n1244), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1238), .B1(new_n744), .B2(new_n1252), .C1(new_n917), .C2(new_n792), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1237), .B(new_n1253), .C1(new_n1161), .C2(new_n737), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n737), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1253), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT122), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1236), .A2(new_n1258), .ZN(G381));
  OR4_X1    g1059(.A1(G396), .A2(G387), .A3(G384), .A4(G393), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1198), .A2(new_n1223), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT57), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1228), .A2(new_n1229), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n700), .B1(new_n1263), .B2(new_n1231), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1262), .B1(new_n1226), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1261), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1171), .A2(new_n699), .A3(new_n1173), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1268), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G390), .A2(new_n1260), .A3(G381), .A4(new_n1270), .ZN(G407));
  NOR2_X1   g1071(.A1(new_n671), .A2(G343), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT123), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(new_n1270), .C2(new_n1274), .ZN(G409));
  XNOR2_X1  g1075(.A(G393), .B(G396), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1276), .A2(new_n1083), .A3(new_n1080), .A4(new_n1104), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G393), .B(new_n809), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G387), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1279), .A3(new_n1039), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1161), .A2(KEYINPUT60), .A3(new_n1163), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n699), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1258), .B(G384), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1288), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n699), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1293), .A2(KEYINPUT124), .A3(G384), .A4(new_n1258), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1258), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1295));
  INV_X1    g1095(.A(G384), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1291), .A2(new_n1294), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G2897), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1274), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1272), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1291), .A2(new_n1297), .A3(new_n1294), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1231), .A2(new_n1234), .A3(new_n1197), .A4(new_n1195), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1198), .A3(new_n1223), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1269), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT115), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1268), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1175), .A2(KEYINPUT115), .A3(new_n1171), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1309), .B1(G375), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1306), .B1(new_n1315), .B2(new_n1274), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1284), .B1(new_n1316), .B2(KEYINPUT61), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1267), .A2(G378), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1273), .B1(new_n1319), .B2(new_n1309), .ZN(new_n1320));
  OAI211_X1 g1120(.A(KEYINPUT127), .B(new_n1318), .C1(new_n1320), .C2(new_n1306), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1298), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1315), .A2(new_n1302), .A3(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1298), .A2(new_n1323), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1323), .A2(new_n1325), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1283), .B1(new_n1322), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1298), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1315), .A2(new_n1274), .A3(new_n1331), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1277), .A2(new_n1279), .A3(new_n1039), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1039), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1333), .A2(new_n1334), .A3(KEYINPUT61), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1272), .B1(new_n1319), .B2(new_n1309), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1332), .B(new_n1335), .C1(new_n1336), .C2(new_n1306), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1339), .B1(new_n1336), .B2(new_n1324), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1329), .B1(new_n1337), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1281), .A2(new_n1318), .A3(new_n1282), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1315), .A2(new_n1302), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1306), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1325), .A2(new_n1338), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(KEYINPUT126), .A4(new_n1332), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1341), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1328), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1269), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1319), .A2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1283), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1324), .ZN(G402));
endmodule


