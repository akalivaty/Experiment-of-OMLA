//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT86), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n210), .A2(new_n212), .B1(KEYINPUT2), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n213), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT82), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n213), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n213), .ZN(new_n224));
  XNOR2_X1  g023(.A(G141gat), .B(G148gat), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT82), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT78), .B(G218gat), .Z(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT29), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n228), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(new_n232), .B2(new_n233), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n223), .B2(new_n227), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(KEYINPUT29), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n208), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n223), .A2(new_n227), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n243), .B2(new_n244), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n206), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n238), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n246), .A2(KEYINPUT29), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(G22gat), .B1(new_n248), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n205), .B1(new_n259), .B2(KEYINPUT88), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n249), .B1(new_n251), .B2(new_n240), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n255), .A2(new_n256), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n207), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n228), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n247), .A3(new_n254), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n264), .A2(new_n267), .A3(KEYINPUT89), .A4(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(G22gat), .C1(new_n248), .C2(new_n258), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n268), .A3(KEYINPUT87), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(G22gat), .C1(new_n248), .C2(new_n258), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n205), .ZN(new_n279));
  OAI22_X1  g078(.A1(new_n261), .A2(new_n274), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT73), .B(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT1), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  INV_X1    g085(.A(G127gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(G134gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G127gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(new_n287), .A3(G134gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n287), .B2(G134gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n289), .A2(G127gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(KEYINPUT72), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G113gat), .A2(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n292), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(G190gat), .B1(new_n311), .B2(KEYINPUT27), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT26), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT69), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n312), .A2(KEYINPUT68), .A3(new_n309), .A4(new_n313), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n315), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT25), .B1(new_n320), .B2(KEYINPUT23), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n325), .A2(KEYINPUT67), .A3(KEYINPUT24), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n340), .A2(G169gat), .A3(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n323), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n323), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n332), .A2(new_n338), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n347), .A3(new_n323), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT64), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT64), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n311), .A3(new_n306), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(new_n325), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n348), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n346), .B1(new_n359), .B2(KEYINPUT25), .ZN(new_n360));
  INV_X1    g159(.A(new_n326), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n308), .A2(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n342), .B1(new_n318), .B2(KEYINPUT26), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n333), .B1(new_n364), .B2(new_n322), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(KEYINPUT70), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n304), .A2(new_n329), .A3(new_n360), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT74), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n344), .A2(new_n347), .A3(new_n323), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n325), .A2(new_n357), .ZN(new_n370));
  INV_X1    g169(.A(new_n356), .ZN(new_n371));
  NOR3_X1   g170(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n350), .A2(new_n352), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(new_n346), .B1(new_n327), .B2(new_n328), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n304), .A4(new_n366), .ZN(new_n380));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n329), .A2(new_n360), .A3(new_n366), .ZN(new_n382));
  INV_X1    g181(.A(new_n304), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n380), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n281), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n390), .A2(new_n386), .A3(KEYINPUT75), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n380), .A3(new_n384), .ZN(new_n393));
  INV_X1    g192(.A(new_n381), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT33), .B1(new_n393), .B2(new_n394), .ZN(new_n396));
  XOR2_X1   g195(.A(G15gat), .B(G43gat), .Z(new_n397));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n395), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  AOI221_X4 g200(.A(new_n392), .B1(KEYINPUT33), .B2(new_n399), .C1(new_n393), .C2(new_n394), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n389), .A2(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n395), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n393), .A2(new_n394), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n407), .A3(new_n399), .ZN(new_n408));
  INV_X1    g207(.A(new_n402), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n390), .A2(new_n386), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n280), .A2(new_n403), .A3(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G1gat), .B(G29gat), .Z(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(new_n303), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n299), .B2(new_n300), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n228), .B1(new_n421), .B2(new_n292), .ZN(new_n422));
  INV_X1    g221(.A(new_n300), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT71), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT72), .B1(new_n424), .B2(new_n294), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n303), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n292), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n249), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n419), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n246), .B1(KEYINPUT3), .B2(new_n228), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n434), .B2(new_n383), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n304), .A2(new_n436), .A3(new_n249), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n304), .A2(KEYINPUT84), .A3(new_n436), .A4(new_n249), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n433), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n437), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n435), .A2(new_n444), .A3(new_n419), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n418), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n435), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n432), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n417), .A3(new_n445), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT6), .B(new_n418), .C1(new_n443), .C2(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n377), .A2(new_n346), .B1(new_n365), .B2(new_n363), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n341), .A2(new_n339), .A3(new_n342), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT66), .B1(new_n344), .B2(new_n323), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n347), .B(KEYINPUT25), .C1(new_n337), .C2(new_n325), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n375), .A2(new_n376), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n327), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT79), .B(new_n459), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n382), .B2(new_n250), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n245), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G64gat), .B(G92gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n472), .B(new_n473), .Z(new_n474));
  AOI21_X1  g273(.A(KEYINPUT29), .B1(new_n360), .B2(new_n327), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n459), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n250), .B1(new_n466), .B2(new_n467), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n457), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n382), .A2(new_n459), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n471), .B(new_n474), .C1(new_n481), .C2(new_n245), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n477), .A3(new_n457), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT80), .B1(new_n475), .B2(new_n459), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n457), .B1(new_n378), .B2(new_n366), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n255), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n471), .A4(new_n474), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n483), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n474), .B1(new_n489), .B2(new_n471), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n458), .A2(new_n468), .ZN(new_n494));
  INV_X1    g293(.A(new_n470), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n255), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n457), .B1(new_n456), .B2(KEYINPUT29), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n480), .A3(KEYINPUT80), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n245), .B1(new_n498), .B2(new_n485), .ZN(new_n499));
  INV_X1    g298(.A(new_n474), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n493), .B1(new_n501), .B2(KEYINPUT30), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n454), .A2(new_n492), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT35), .B1(new_n412), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n505));
  AND4_X1   g304(.A1(new_n454), .A2(new_n492), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n387), .A2(new_n388), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n401), .B2(new_n402), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n411), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n510));
  INV_X1    g309(.A(new_n279), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n510), .A2(new_n260), .B1(new_n275), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n408), .A2(new_n409), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n387), .A2(new_n281), .A3(new_n388), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT75), .B1(new_n390), .B2(new_n386), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT76), .B1(new_n520), .B2(new_n411), .ZN(new_n521));
  AND4_X1   g320(.A1(KEYINPUT76), .A2(new_n403), .A3(KEYINPUT36), .A4(new_n411), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n509), .B2(new_n515), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT77), .B(KEYINPUT36), .C1(new_n508), .C2(new_n411), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n521), .A2(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n441), .A2(new_n437), .B1(new_n434), .B2(new_n383), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT39), .B1(new_n528), .B2(new_n430), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n422), .A2(new_n428), .A3(new_n430), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n434), .A2(new_n383), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n436), .B1(new_n304), .B2(new_n249), .ZN(new_n535));
  AND4_X1   g334(.A1(new_n436), .A2(new_n426), .A3(new_n427), .A4(new_n249), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT39), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n431), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n417), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n527), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n447), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n430), .B1(new_n444), .B2(new_n534), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n418), .B1(new_n543), .B2(new_n538), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(KEYINPUT40), .C1(new_n532), .C2(new_n529), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n529), .A2(new_n532), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n544), .A3(new_n548), .A4(KEYINPUT40), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n542), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n492), .A2(new_n502), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n512), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n452), .A2(new_n453), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n474), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n493), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n481), .A2(new_n255), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n255), .B1(new_n469), .B2(new_n470), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT37), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n554), .B1(new_n489), .B2(new_n471), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT38), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n483), .A2(new_n491), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n553), .A2(new_n562), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n552), .A2(new_n566), .B1(new_n503), .B2(new_n512), .ZN(new_n567));
  AOI221_X4 g366(.A(new_n202), .B1(new_n504), .B2(new_n514), .C1(new_n526), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n526), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n514), .A2(new_n504), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT93), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G8gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT94), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT16), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(G1gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n577), .B2(KEYINPUT95), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(G1gat), .B2(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI221_X1 g379(.A(new_n577), .B1(KEYINPUT95), .B2(new_n573), .C1(G1gat), .C2(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n582), .B1(KEYINPUT21), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT98), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT99), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n592), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G36gat), .ZN(new_n602));
  AND2_X1   g401(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G29gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n610));
  XNOR2_X1  g409(.A(G43gat), .B(G50gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT8), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(KEYINPUT101), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(G99gat), .A3(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n617), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT100), .B(new_n623), .C1(new_n620), .C2(new_n621), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT100), .B1(new_n620), .B2(new_n621), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(G85gat), .A3(G92gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT7), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G99gat), .B(G106gat), .Z(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n636), .B2(new_n613), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G190gat), .B(G218gat), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n641), .A3(new_n637), .ZN(new_n642));
  XOR2_X1   g441(.A(G134gat), .B(G162gat), .Z(new_n643));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT103), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n638), .A2(new_n639), .B1(KEYINPUT102), .B2(new_n646), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n642), .A3(new_n650), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n601), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n587), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  INV_X1    g456(.A(new_n587), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n636), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n659), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(G120gat), .B(G148gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n664), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n662), .B2(new_n663), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT105), .B(new_n666), .C1(new_n660), .C2(new_n661), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n667), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n671), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n655), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n652), .A2(new_n654), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n592), .B(new_n599), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n679), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n582), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n614), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G229gat), .A2(G233gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT96), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n582), .A2(new_n613), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT18), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n689), .A2(KEYINPUT18), .A3(new_n691), .A4(new_n692), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n582), .B(new_n613), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n691), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(G113gat), .B(G141gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G197gat), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT11), .B(G169gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT12), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n706), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n695), .A2(new_n708), .A3(new_n696), .A4(new_n700), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n687), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n572), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n553), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g513(.A1(new_n572), .A2(new_n551), .A3(new_n711), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n576), .A2(new_n573), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n718), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n715), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(G1325gat));
  AND2_X1   g523(.A1(new_n508), .A2(new_n411), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT77), .B1(new_n725), .B2(KEYINPUT36), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n509), .A2(new_n523), .A3(new_n515), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n403), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT76), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n520), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n726), .A2(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n712), .A2(G15gat), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(G15gat), .B1(new_n712), .B2(new_n725), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(G1326gat));
  NAND2_X1  g536(.A1(new_n712), .A2(new_n512), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT43), .B(G22gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  NAND2_X1  g539(.A1(new_n503), .A2(new_n512), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n492), .A2(new_n502), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n546), .A2(new_n549), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n541), .A2(new_n447), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n280), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n483), .B(new_n491), .C1(new_n556), .C2(new_n561), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n500), .B1(new_n496), .B2(new_n499), .ZN(new_n748));
  INV_X1    g547(.A(new_n555), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n563), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n557), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n747), .A2(new_n752), .A3(new_n454), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n741), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n570), .B1(new_n732), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n202), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n569), .A2(KEYINPUT93), .A3(new_n570), .ZN(new_n757));
  INV_X1    g556(.A(new_n710), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n601), .A3(new_n680), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n756), .A2(new_n757), .A3(new_n682), .A4(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(G29gat), .A3(new_n454), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT45), .Z(new_n762));
  NAND3_X1  g561(.A1(new_n756), .A2(new_n757), .A3(new_n682), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n514), .A2(new_n504), .A3(KEYINPUT109), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT109), .B1(new_n514), .B2(new_n504), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n569), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(new_n768), .A3(new_n682), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n759), .ZN(new_n771));
  OAI21_X1  g570(.A(G29gat), .B1(new_n771), .B2(new_n454), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n762), .A2(new_n772), .ZN(G1328gat));
  OAI21_X1  g572(.A(G36gat), .B1(new_n771), .B2(new_n742), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n760), .A2(G36gat), .A3(new_n742), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1329gat));
  AND4_X1   g576(.A1(G43gat), .A2(new_n770), .A3(new_n732), .A4(new_n759), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n509), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(G43gat), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT47), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1330gat));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n768), .B1(new_n572), .B2(new_n682), .ZN(new_n786));
  INV_X1    g585(.A(new_n769), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n512), .B(new_n759), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n788), .B2(G50gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n760), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n280), .A2(G50gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n760), .B2(new_n790), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT112), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n572), .A2(KEYINPUT111), .A3(new_n682), .A4(new_n759), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n760), .A2(new_n790), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n788), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n795), .A2(new_n796), .A3(new_n792), .ZN(new_n802));
  INV_X1    g601(.A(new_n785), .ZN(new_n803));
  INV_X1    g602(.A(new_n759), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n280), .B(new_n804), .C1(new_n764), .C2(new_n769), .ZN(new_n805));
  INV_X1    g604(.A(G50gat), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n802), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n800), .A2(new_n801), .B1(KEYINPUT48), .B2(new_n807), .ZN(G1331gat));
  AND4_X1   g607(.A1(new_n684), .A2(new_n767), .A3(new_n680), .A4(new_n758), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n553), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n551), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT49), .B(G64gat), .Z(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(G1333gat));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n732), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n509), .A2(G71gat), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n816), .A2(G71gat), .B1(new_n809), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g618(.A1(new_n809), .A2(new_n512), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g620(.A1(new_n710), .A2(new_n601), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n680), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n764), .B2(new_n769), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825), .B2(new_n454), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n767), .A2(new_n682), .A3(new_n822), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n679), .A2(new_n454), .A3(G85gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n826), .A2(new_n834), .ZN(G1336gat));
  NOR3_X1   g634(.A1(new_n742), .A2(G92gat), .A3(new_n679), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n829), .B2(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n824), .A2(new_n551), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(G92gat), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n841), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n838), .C1(new_n839), .C2(G92gat), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(new_n844), .ZN(G1337gat));
  OAI21_X1  g644(.A(G99gat), .B1(new_n825), .B2(new_n526), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n509), .A2(new_n679), .A3(G99gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1338gat));
  INV_X1    g648(.A(G106gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n824), .B2(new_n512), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n679), .A2(new_n280), .A3(G106gat), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n831), .A2(new_n852), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1339gat));
  INV_X1    g655(.A(new_n675), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n662), .A2(new_n674), .A3(new_n663), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n662), .B2(new_n663), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n660), .A2(new_n666), .A3(new_n661), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n671), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n860), .A2(KEYINPUT55), .A3(new_n863), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n710), .A3(new_n672), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n697), .A2(new_n699), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n691), .B1(new_n689), .B2(new_n692), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n705), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n709), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n679), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n682), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n682), .A2(new_n709), .A3(new_n871), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n672), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT55), .B1(new_n860), .B2(new_n863), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n683), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n684), .A2(new_n758), .A3(new_n679), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n454), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n412), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n742), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n282), .A3(new_n710), .ZN(new_n886));
  INV_X1    g685(.A(new_n513), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n880), .B2(new_n881), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n742), .A2(new_n553), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G113gat), .B1(new_n892), .B2(new_n758), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n886), .A2(new_n893), .ZN(G1340gat));
  AOI21_X1  g693(.A(G120gat), .B1(new_n885), .B2(new_n680), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n679), .A2(new_n283), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n891), .B2(new_n896), .ZN(G1341gat));
  NAND3_X1  g696(.A1(new_n885), .A2(new_n287), .A3(new_n601), .ZN(new_n898));
  OAI21_X1  g697(.A(G127gat), .B1(new_n892), .B2(new_n683), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1342gat));
  INV_X1    g699(.A(new_n682), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n551), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n884), .A2(new_n289), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT115), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(KEYINPUT115), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n682), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n908), .B2(G134gat), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n906), .B(new_n907), .C1(new_n909), .C2(new_n903), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n732), .A2(new_n890), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n280), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n881), .ZN(new_n915));
  XOR2_X1   g714(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n916));
  AOI22_X1  g715(.A1(new_n864), .A2(new_n916), .B1(new_n707), .B2(new_n709), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n867), .A2(new_n672), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n873), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n866), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n919), .A2(new_n682), .B1(new_n920), .B2(new_n876), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n683), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(KEYINPUT117), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n924), .A3(new_n683), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n914), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n880), .A2(new_n881), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n512), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n911), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G141gat), .B1(new_n929), .B2(new_n758), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n732), .A2(new_n280), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n882), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(new_n742), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n209), .A3(new_n710), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT58), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n930), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1344gat));
  OR3_X1    g738(.A1(new_n929), .A2(KEYINPUT59), .A3(new_n679), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n911), .A2(new_n680), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n921), .A2(new_n683), .B1(new_n687), .B2(new_n758), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n512), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n687), .A2(new_n758), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n922), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n912), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n913), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n933), .B2(new_n680), .ZN(new_n952));
  OAI221_X1 g751(.A(new_n940), .B1(new_n949), .B2(new_n950), .C1(new_n952), .C2(G148gat), .ZN(G1345gat));
  NOR2_X1   g752(.A1(new_n683), .A2(new_n218), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT119), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n929), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(G155gat), .B1(new_n933), .B2(new_n601), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n929), .B2(new_n901), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n932), .A2(new_n219), .A3(new_n902), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n742), .A2(new_n553), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n927), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n883), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT120), .Z(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n710), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n963), .B(KEYINPUT121), .Z(new_n968));
  NOR2_X1   g767(.A1(new_n889), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n758), .A2(new_n316), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n967), .A2(new_n316), .B1(new_n969), .B2(new_n970), .ZN(G1348gat));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n317), .A3(new_n680), .ZN(new_n972));
  INV_X1    g771(.A(new_n969), .ZN(new_n973));
  OAI21_X1  g772(.A(G176gat), .B1(new_n973), .B2(new_n679), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1349gat));
  INV_X1    g774(.A(new_n968), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n927), .A2(new_n513), .A3(new_n601), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT122), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n888), .A2(new_n979), .A3(new_n601), .A4(new_n976), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(G183gat), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(new_n313), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n964), .A2(new_n883), .A3(new_n601), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT124), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n987), .A2(KEYINPUT123), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n981), .A2(new_n989), .A3(new_n984), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n986), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(G1350gat));
  NAND3_X1  g792(.A1(new_n966), .A2(new_n306), .A3(new_n682), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n306), .B1(new_n969), .B2(new_n682), .ZN(new_n995));
  XNOR2_X1  g794(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(G1351gat));
  AND2_X1   g797(.A1(new_n964), .A2(new_n931), .ZN(new_n999));
  AOI21_X1  g798(.A(G197gat), .B1(new_n999), .B2(new_n710), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n968), .A2(new_n732), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT126), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1002), .B1(new_n947), .B2(new_n948), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n710), .A2(G197gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(G1352gat));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  INV_X1    g805(.A(G204gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n1003), .B2(new_n680), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n964), .A2(new_n1007), .A3(new_n680), .A4(new_n931), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1009), .B(KEYINPUT62), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(new_n1002), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n922), .A2(new_n945), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n280), .B1(new_n1013), .B2(KEYINPUT118), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n942), .A2(new_n943), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT57), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(new_n948), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n680), .B(new_n1012), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(G204gat), .ZN(new_n1019));
  XOR2_X1   g818(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1020));
  NAND3_X1  g819(.A1(new_n1019), .A2(new_n1020), .A3(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1011), .A2(new_n1021), .ZN(G1353gat));
  NAND3_X1  g821(.A1(new_n999), .A2(new_n231), .A3(new_n601), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n601), .B(new_n1012), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  AOI21_X1  g826(.A(G218gat), .B1(new_n999), .B2(new_n682), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n901), .A2(new_n230), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1028), .B1(new_n1003), .B2(new_n1029), .ZN(G1355gat));
endmodule


