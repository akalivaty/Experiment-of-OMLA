//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(G1gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210));
  AOI21_X1  g009(.A(G8gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n211), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n220), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G43gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT86), .B(G43gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G50gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(G43gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(KEYINPUT15), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n221), .A2(new_n229), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n215), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT13), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(new_n215), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n231), .A2(KEYINPUT17), .A3(new_n232), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n241), .A2(new_n215), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(KEYINPUT17), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(new_n235), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n238), .B1(new_n245), .B2(KEYINPUT18), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n207), .B1(new_n246), .B2(KEYINPUT88), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n246), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n249), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g057(.A1(G113gat), .A2(G120gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n258), .A4(new_n259), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G127gat), .ZN(new_n263));
  INV_X1    g062(.A(G127gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G134gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n254), .A2(new_n260), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n260), .A2(new_n254), .A3(new_n266), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT74), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n254), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n260), .A2(new_n254), .A3(new_n266), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n277));
  NOR2_X1   g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT24), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n204), .A2(new_n284), .A3(KEYINPUT23), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n277), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT66), .B(new_n277), .C1(new_n283), .C2(new_n289), .ZN(new_n293));
  INV_X1    g092(.A(new_n289), .ZN(new_n294));
  OR2_X1    g093(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n280), .A2(new_n282), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n294), .B(KEYINPUT25), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n292), .A2(new_n293), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n204), .A2(new_n284), .A3(KEYINPUT71), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n302), .A2(KEYINPUT26), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n279), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT27), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n308), .A3(KEYINPUT27), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n310), .A2(new_n312), .A3(new_n295), .A4(new_n296), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n307), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT67), .B(G190gat), .Z(new_n318));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT28), .A4(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n295), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n306), .B1(new_n317), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n276), .B1(new_n301), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n317), .ZN(new_n330));
  INV_X1    g129(.A(new_n306), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n292), .A2(new_n293), .A3(new_n300), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n269), .A4(new_n275), .ZN(new_n334));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT64), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT33), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT75), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  AOI211_X1 g145(.A(new_n346), .B(new_n343), .C1(new_n337), .C2(new_n339), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n344), .B2(KEYINPUT33), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n337), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n334), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT34), .ZN(new_n352));
  INV_X1    g151(.A(new_n336), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n329), .A2(new_n334), .B1(G227gat), .B2(G233gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n350), .B(new_n354), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n358), .B(new_n359), .C1(new_n345), .C2(new_n347), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G211gat), .B(G218gat), .Z(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT77), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n364), .B1(KEYINPUT22), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n363), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G226gat), .ZN(new_n370));
  INV_X1    g169(.A(G233gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n332), .A2(new_n333), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n370), .B(new_n371), .C1(new_n332), .C2(new_n333), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n372), .ZN(new_n378));
  INV_X1    g177(.A(new_n369), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n332), .B2(new_n333), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n378), .B(new_n379), .C1(new_n372), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G64gat), .ZN(new_n383));
  INV_X1    g182(.A(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(KEYINPUT30), .Z(new_n386));
  AND3_X1   g185(.A1(new_n377), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(KEYINPUT30), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n377), .B2(new_n381), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(G141gat), .ZN(new_n392));
  INV_X1    g191(.A(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395));
  AND2_X1   g194(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n396));
  NOR2_X1   g195(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n394), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n404));
  INV_X1    g203(.A(G155gat), .ZN(new_n405));
  INV_X1    g204(.A(G162gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  AND2_X1   g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(KEYINPUT79), .A3(new_n395), .ZN(new_n412));
  AOI221_X4 g211(.A(new_n403), .B1(new_n399), .B2(new_n407), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n412), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n407), .A2(new_n399), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT80), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n402), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n272), .A2(new_n274), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n267), .A2(new_n268), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n402), .C1(new_n416), .C2(new_n413), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n391), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  INV_X1    g225(.A(new_n402), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n409), .A2(new_n410), .A3(new_n408), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT79), .B1(new_n394), .B2(new_n395), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n415), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n403), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n414), .A2(KEYINPUT80), .A3(new_n415), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n426), .B1(new_n276), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n418), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n417), .A2(KEYINPUT3), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n423), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n425), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n421), .A2(KEYINPUT4), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n276), .A2(new_n426), .A3(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n420), .B1(new_n417), .B2(KEYINPUT3), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n433), .A2(new_n437), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n444), .A2(new_n423), .A3(new_n447), .A4(new_n391), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT0), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G57gat), .ZN(new_n452));
  INV_X1    g251(.A(G85gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n448), .A3(new_n454), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n390), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n350), .B1(new_n345), .B2(new_n347), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n354), .B1(new_n352), .B2(new_n355), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G78gat), .B(G106gat), .Z(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n379), .B1(new_n446), .B2(new_n374), .ZN(new_n469));
  INV_X1    g268(.A(new_n362), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n368), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT29), .B1(new_n368), .B2(new_n470), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT3), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n433), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n369), .B1(new_n439), .B2(KEYINPUT29), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n437), .B1(new_n369), .B2(KEYINPUT29), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n468), .B1(new_n477), .B2(new_n417), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  INV_X1    g280(.A(G22gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n467), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n475), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n475), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G22gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n475), .B2(new_n479), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n480), .A2(KEYINPUT82), .A3(new_n482), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n467), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n486), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n361), .A2(new_n461), .A3(new_n464), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n358), .B1(new_n345), .B2(new_n347), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n464), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n390), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n459), .B2(new_n460), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n494), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n464), .A2(new_n498), .A3(KEYINPUT36), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n357), .A2(new_n360), .B1(new_n462), .B2(new_n463), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(KEYINPUT36), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n461), .A2(new_n494), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n454), .B1(new_n441), .B2(new_n448), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n509), .A2(new_n387), .A3(new_n389), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT39), .B1(new_n422), .B2(new_n424), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n444), .A2(new_n447), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(new_n424), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n442), .A2(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n423), .A2(KEYINPUT39), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n454), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n511), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n512), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n423), .B2(new_n515), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n455), .B1(new_n513), .B2(new_n516), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT40), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT84), .A4(KEYINPUT40), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n519), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n459), .A2(new_n460), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT37), .B1(new_n377), .B2(new_n381), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT37), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n385), .A2(new_n533), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n377), .A2(KEYINPUT37), .A3(new_n381), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n529), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n377), .A2(new_n381), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n385), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n527), .B(new_n494), .C1(new_n528), .C2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n507), .A2(new_n508), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n253), .B1(new_n504), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(G71gat), .ZN(new_n546));
  INV_X1    g345(.A(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G64gat), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(KEYINPUT90), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(KEYINPUT90), .B2(new_n554), .ZN(new_n556));
  INV_X1    g355(.A(new_n549), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n551), .B(new_n556), .C1(KEYINPUT9), .C2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT92), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT9), .B1(new_n554), .B2(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n557), .B1(new_n561), .B2(new_n548), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n560), .B(new_n562), .C1(new_n561), .C2(new_n548), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n453), .B2(new_n384), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G99gat), .B(G106gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n559), .A2(new_n563), .ZN(new_n574));
  INV_X1    g373(.A(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT98), .A3(new_n571), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n577), .A2(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n545), .B(new_n573), .C1(new_n582), .C2(KEYINPUT10), .ZN(new_n583));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G176gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(G204gat), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n577), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n581), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n545), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(KEYINPUT99), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(KEYINPUT99), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n583), .B(new_n586), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n583), .A2(new_n591), .ZN(new_n595));
  INV_X1    g394(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT100), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  AOI211_X1 g397(.A(new_n598), .B(new_n586), .C1(new_n583), .C2(new_n591), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n215), .B1(new_n574), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G183gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n574), .A2(new_n601), .ZN(new_n608));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n365), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n243), .A2(new_n241), .A3(new_n575), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n233), .A2(new_n571), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT93), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT96), .Z(new_n626));
  AOI21_X1  g425(.A(new_n619), .B1(new_n626), .B2(KEYINPUT95), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n622), .A2(new_n624), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT94), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n600), .A2(new_n615), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n544), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n528), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n390), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT16), .B(G8gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(G8gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n635), .B2(new_n507), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n361), .A2(new_n464), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(G15gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n635), .B2(new_n649), .ZN(G1326gat));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n494), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT43), .B(G22gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT101), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n504), .A2(new_n543), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n633), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n541), .A2(new_n528), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n525), .A2(new_n526), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n390), .A2(new_n456), .A3(new_n519), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n494), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI22_X1  g462(.A1(new_n660), .A2(new_n663), .B1(new_n461), .B2(new_n494), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n464), .A2(KEYINPUT36), .A3(new_n498), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n648), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n659), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n507), .A2(new_n542), .A3(KEYINPUT102), .A4(new_n508), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT103), .B1(new_n670), .B2(new_n504), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n672), .B(new_n503), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n633), .A2(new_n656), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n658), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n600), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n615), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n253), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n655), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT104), .B(new_n680), .C1(new_n683), .C2(new_n658), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n528), .ZN(new_n686));
  INV_X1    g485(.A(new_n679), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n633), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(new_n216), .A3(new_n637), .A4(new_n544), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(G1328gat));
  OAI21_X1  g491(.A(G36gat), .B1(new_n685), .B2(new_n500), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n689), .A2(new_n217), .A3(new_n390), .A4(new_n544), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT46), .Z(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n689), .A2(new_n506), .A3(new_n224), .A4(new_n544), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n677), .A2(new_n507), .A3(new_n681), .ZN(new_n699));
  INV_X1    g498(.A(new_n224), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT47), .ZN(new_n701));
  OAI221_X1 g500(.A(new_n697), .B1(new_n698), .B2(KEYINPUT47), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n697), .A2(new_n698), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n682), .A2(new_n667), .A3(new_n684), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n700), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n705), .B2(KEYINPUT47), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n702), .B(KEYINPUT106), .C1(new_n705), .C2(KEYINPUT47), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  INV_X1    g509(.A(new_n494), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n222), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT107), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n689), .A2(new_n544), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n677), .A2(new_n494), .A3(new_n681), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n222), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n682), .A2(new_n711), .A3(new_n684), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n714), .B1(new_n719), .B2(G50gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g520(.A1(new_n671), .A2(new_n673), .ZN(new_n722));
  INV_X1    g521(.A(new_n633), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n253), .A3(new_n614), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n722), .A2(new_n678), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n637), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  INV_X1    g526(.A(new_n725), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n500), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  OAI21_X1  g532(.A(new_n546), .B1(new_n728), .B2(new_n648), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n725), .A2(G71gat), .A3(new_n667), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n725), .A2(new_n711), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n614), .A2(new_n742), .A3(new_n252), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT109), .B1(new_n615), .B2(new_n253), .ZN(new_n744));
  OAI221_X1 g543(.A(new_n600), .B1(new_n743), .B2(new_n744), .C1(new_n683), .C2(new_n658), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n528), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n633), .B1(new_n744), .B2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n503), .B1(new_n668), .B2(new_n669), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n678), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n453), .A3(new_n637), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n753), .ZN(G1336gat));
  OAI21_X1  g553(.A(G92gat), .B1(new_n745), .B2(new_n500), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n500), .A2(G92gat), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n752), .A2(KEYINPUT111), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n752), .B2(new_n757), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n755), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n752), .A2(new_n757), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n757), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n755), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n765), .B2(new_n756), .ZN(G1337gat));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n745), .A2(new_n767), .A3(new_n507), .ZN(new_n768));
  AOI21_X1  g567(.A(G99gat), .B1(new_n752), .B2(new_n506), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1338gat));
  OAI21_X1  g569(.A(G106gat), .B1(new_n745), .B2(new_n494), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT53), .B1(new_n771), .B2(KEYINPUT113), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n750), .A2(new_n751), .ZN(new_n773));
  OR3_X1    g572(.A1(new_n678), .A2(G106gat), .A3(new_n494), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT112), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n772), .B(new_n776), .Z(G1339gat));
  NAND2_X1  g576(.A1(new_n506), .A2(new_n494), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n248), .A2(new_n246), .A3(new_n207), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n234), .A2(new_n237), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT114), .Z(new_n781));
  NOR2_X1   g580(.A1(new_n244), .A2(new_n235), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n206), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n600), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT10), .B1(new_n587), .B2(new_n588), .ZN(new_n786));
  INV_X1    g585(.A(new_n573), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n590), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n583), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n596), .B1(new_n583), .B2(KEYINPUT54), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n583), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n786), .A2(new_n787), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n545), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n792), .A2(new_n795), .A3(KEYINPUT55), .A4(new_n596), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n791), .A2(new_n252), .A3(new_n594), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n633), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n791), .A2(new_n594), .A3(new_n796), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n633), .A2(new_n779), .A3(new_n783), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n615), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n724), .A2(new_n600), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n778), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n528), .A2(new_n390), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(new_n255), .A3(new_n253), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n528), .B1(new_n802), .B2(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n499), .A2(new_n494), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n390), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n252), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n807), .B1(new_n255), .B2(new_n813), .ZN(G1340gat));
  NOR3_X1   g613(.A1(new_n806), .A2(new_n256), .A3(new_n678), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n600), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n256), .B2(new_n816), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n806), .B2(new_n615), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n614), .A2(new_n264), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n811), .B2(new_n819), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n723), .A2(G134gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n808), .A2(new_n810), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n806), .B2(new_n723), .ZN(new_n828));
  AOI211_X1 g627(.A(KEYINPUT116), .B(new_n825), .C1(new_n824), .C2(new_n826), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n822), .B(new_n823), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(KEYINPUT56), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n832), .ZN(G1343gat));
  AOI21_X1  g632(.A(new_n494), .B1(new_n802), .B2(new_n803), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT57), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n507), .A2(new_n805), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G141gat), .B1(new_n838), .B2(new_n253), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n507), .A2(new_n711), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n390), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n808), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(G141gat), .A3(new_n253), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n802), .A2(new_n803), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n711), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n849), .A2(new_n837), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n392), .B1(new_n852), .B2(new_n252), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT58), .B1(new_n853), .B2(new_n844), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n854), .ZN(G1344gat));
  INV_X1    g654(.A(new_n843), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n393), .A3(new_n600), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n836), .B(KEYINPUT117), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n849), .A2(new_n600), .A3(new_n851), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n393), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n835), .A2(KEYINPUT118), .A3(new_n600), .A4(new_n859), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT59), .B(new_n393), .C1(new_n852), .C2(new_n600), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(G1345gat));
  OAI21_X1  g665(.A(G155gat), .B1(new_n838), .B2(new_n615), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n856), .A2(new_n405), .A3(new_n614), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n838), .B2(new_n723), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n856), .A2(new_n406), .A3(new_n633), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n637), .B1(new_n802), .B2(new_n803), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n809), .A2(new_n500), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n252), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n637), .A2(new_n500), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n804), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n253), .A2(new_n204), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1348gat));
  NOR2_X1   g680(.A1(new_n678), .A2(new_n284), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n284), .B1(new_n875), .B2(new_n678), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(KEYINPUT119), .A3(new_n882), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1349gat));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n320), .A3(new_n614), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n804), .A2(new_n614), .A3(new_n878), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G183gat), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n892), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(KEYINPUT60), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(G1350gat));
  NAND2_X1  g702(.A1(new_n879), .A2(new_n633), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G190gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n875), .A2(new_n297), .A3(new_n723), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT122), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n841), .A2(new_n500), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n873), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(KEYINPUT123), .B(G197gat), .Z(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n252), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n849), .A2(new_n851), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n507), .A2(new_n878), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT124), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n914), .A2(new_n253), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(new_n912), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n835), .A2(new_n600), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n919), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n678), .A2(G204gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n925));
  OAI221_X1 g724(.A(new_n920), .B1(KEYINPUT62), .B2(new_n922), .C1(new_n924), .C2(new_n925), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n365), .A3(new_n614), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT126), .Z(new_n928));
  NAND3_X1  g727(.A1(new_n614), .A2(new_n507), .A3(new_n878), .ZN(new_n929));
  OAI21_X1  g728(.A(G211gat), .B1(new_n914), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT63), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT63), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n911), .B2(new_n633), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n916), .A2(new_n366), .A3(new_n723), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n936), .A2(new_n937), .B1(new_n835), .B2(new_n938), .ZN(G1355gat));
endmodule


