//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  AND2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(KEYINPUT22), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G148gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(G141gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT79), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n222), .ZN(new_n227));
  AND2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT78), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n220), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n222), .B1(new_n225), .B2(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n224), .A2(new_n231), .B1(new_n237), .B2(new_n238), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n210), .A2(KEYINPUT29), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n204), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n233), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n210), .A2(KEYINPUT85), .A3(KEYINPUT29), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n245), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n204), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n253), .B1(new_n212), .B2(new_n242), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n248), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G22gat), .ZN(new_n261));
  XOR2_X1   g060(.A(G78gat), .B(G106gat), .Z(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  AND4_X1   g063(.A1(KEYINPUT86), .A2(new_n257), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n267), .A2(new_n264), .B1(new_n257), .B2(new_n261), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT71), .ZN(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G183gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(G190gat), .B1(new_n274), .B2(G183gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT28), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G183gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT27), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n283), .A2(new_n277), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n278), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  OR3_X1    g084(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g095(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n296), .A2(new_n297), .B1(new_n289), .B2(new_n290), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n299), .A2(new_n301), .B1(new_n279), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n280), .A2(new_n282), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n301), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n295), .A2(new_n311), .B1(new_n314), .B2(new_n288), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n315), .A3(KEYINPUT25), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n285), .A2(new_n293), .B1(new_n304), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n319));
  OAI21_X1  g118(.A(G134gat), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(G127gat), .A2(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G113gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G120gat), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT1), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT68), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n320), .A4(new_n321), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(new_n335), .A3(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n327), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n304), .A2(new_n316), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n283), .B2(new_n277), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n276), .A2(KEYINPUT28), .A3(new_n277), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n292), .B(new_n291), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n328), .A2(new_n333), .B1(new_n337), .B2(new_n339), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT64), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n273), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n352), .A2(new_n355), .A3(KEYINPUT32), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n352), .B2(KEYINPUT32), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n354), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(KEYINPUT32), .C1(new_n353), .C2(new_n273), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n351), .B1(new_n342), .B2(new_n349), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT34), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n352), .A2(KEYINPUT32), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT70), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n355), .A3(KEYINPUT32), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n360), .B1(new_n370), .B2(new_n354), .ZN(new_n371));
  INV_X1    g170(.A(new_n361), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n365), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n269), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n212), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n379), .B(KEYINPUT74), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n343), .A2(new_n346), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n380), .A2(KEYINPUT29), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n347), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n384), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n317), .A2(new_n380), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n212), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT76), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n396), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n390), .A2(new_n212), .A3(new_n391), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n343), .A2(new_n346), .A3(new_n383), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n383), .B1(new_n343), .B2(new_n346), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n380), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n212), .B1(new_n406), .B2(new_n387), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n402), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n389), .A2(KEYINPUT30), .A3(new_n392), .A4(new_n396), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(KEYINPUT77), .A3(new_n398), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n334), .A2(new_n244), .A3(new_n340), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT4), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n348), .A2(new_n423), .A3(new_n244), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n227), .A2(new_n230), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n219), .A2(new_n220), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n428), .A2(new_n213), .B1(KEYINPUT2), .B2(new_n222), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n221), .ZN(new_n430));
  INV_X1    g229(.A(new_n239), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n341), .A2(new_n432), .A3(new_n240), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n423), .B1(new_n348), .B2(new_n244), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n425), .A2(new_n426), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n341), .A2(new_n245), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n420), .ZN(new_n439));
  INV_X1    g238(.A(new_n426), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n419), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n433), .A2(new_n437), .A3(new_n426), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  AND4_X1   g244(.A1(new_n423), .A2(new_n334), .A3(new_n244), .A4(new_n340), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n434), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n421), .A2(KEYINPUT82), .A3(new_n424), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n443), .B(new_n444), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  INV_X1    g249(.A(new_n444), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT83), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n442), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n446), .A2(new_n434), .A3(new_n445), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT82), .B1(new_n421), .B2(new_n424), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n443), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n457), .A2(new_n458), .B1(new_n436), .B2(new_n441), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n418), .B(KEYINPUT87), .Z(new_n460));
  OAI211_X1 g259(.A(new_n414), .B(new_n453), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n441), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n449), .B2(new_n452), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT35), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n377), .A2(new_n413), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n414), .B(new_n453), .C1(new_n459), .C2(new_n418), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT84), .B(new_n412), .C1(new_n467), .C2(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n457), .A2(new_n458), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n418), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n414), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n469), .B1(new_n473), .B2(new_n413), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n468), .A2(new_n474), .A3(new_n376), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n479));
  INV_X1    g278(.A(new_n363), .ZN(new_n480));
  AOI211_X1 g279(.A(new_n480), .B(new_n374), .C1(new_n359), .C2(new_n361), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n375), .A2(KEYINPUT36), .A3(new_n366), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n389), .A2(new_n392), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n402), .B1(new_n487), .B2(KEYINPUT37), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n389), .B2(new_n392), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n397), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n408), .B1(new_n489), .B2(new_n396), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n390), .A2(new_n378), .A3(new_n391), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(KEYINPUT37), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n212), .B1(new_n385), .B2(new_n388), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n461), .A2(new_n464), .A3(new_n491), .A4(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n433), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n447), .B2(new_n448), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n440), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT88), .B1(new_n439), .B2(new_n440), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n438), .A2(new_n506), .A3(new_n420), .A4(new_n426), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(KEYINPUT39), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n508), .C1(new_n501), .C2(new_n426), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n509), .A3(new_n460), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT40), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n460), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n463), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n512), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n504), .A2(new_n509), .A3(new_n460), .A4(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n513), .A2(new_n412), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n269), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n484), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n265), .A2(new_n268), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n468), .B2(new_n474), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n477), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT11), .B(G169gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT12), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(KEYINPUT96), .C1(G1gat), .C2(new_n532), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT95), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT93), .B(G43gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G50gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(G29gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G36gat), .ZN(new_n545));
  NOR3_X1   g344(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(new_n543), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n546), .B2(KEYINPUT91), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n545), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT15), .A3(new_n542), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n538), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n552), .A2(new_n538), .A3(new_n556), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT17), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n552), .B2(new_n556), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n537), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n559), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n557), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n537), .B(KEYINPUT97), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n558), .A2(new_n559), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n568), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n564), .B(KEYINPUT13), .Z(new_n576));
  AOI22_X1  g375(.A1(new_n569), .A2(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n531), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n577), .A3(new_n531), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT98), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n578), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n525), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT105), .B(G92gat), .Z(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  INV_X1    g393(.A(G99gat), .ZN(new_n595));
  INV_X1    g394(.A(G106gat), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT8), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n561), .B1(new_n565), .B2(new_n557), .ZN(new_n601));
  INV_X1    g400(.A(new_n562), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n573), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n589), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT107), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n607), .B1(new_n560), .B2(new_n562), .ZN(new_n612));
  INV_X1    g411(.A(new_n589), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n566), .A2(new_n600), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT106), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT104), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n611), .B2(new_n616), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n588), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n609), .B(KEYINPUT107), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n615), .B(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n618), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n587), .A3(new_n620), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G57gat), .B(G64gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT100), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G71gat), .B(G78gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G64gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G57gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT101), .B(G57gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(new_n638), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n641), .A3(new_n635), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n567), .B1(KEYINPUT21), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT21), .B1(new_n637), .B2(new_n642), .ZN(new_n647));
  XOR2_X1   g446(.A(G127gat), .B(G155gat), .Z(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n646), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n650), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n645), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n643), .B(new_n600), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n664), .A2(new_n661), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n660), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT109), .Z(new_n671));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n660), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n672), .B2(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n629), .A2(new_n657), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n586), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n473), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n412), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G8gat), .B1(new_n680), .B2(new_n413), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g487(.A(new_n686), .B(new_n688), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n680), .B2(new_n484), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n375), .A2(new_n366), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n680), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n680), .A2(new_n269), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n477), .A2(new_n524), .ZN(new_n699));
  INV_X1    g498(.A(new_n628), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n587), .B1(new_n627), .B2(new_n620), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n520), .B1(new_n523), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(KEYINPUT110), .B(new_n522), .C1(new_n468), .C2(new_n474), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n473), .A2(new_n413), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT84), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n473), .A2(new_n469), .A3(new_n413), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n377), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT35), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n706), .A2(new_n707), .B1(new_n712), .B2(new_n466), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n623), .A2(new_n698), .A3(new_n628), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n704), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n523), .A2(new_n705), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n521), .A3(new_n707), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n477), .ZN(new_n718));
  INV_X1    g517(.A(new_n714), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(KEYINPUT111), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n703), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n676), .A2(new_n657), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n583), .A2(new_n578), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n697), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n525), .B2(new_n629), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT111), .B1(new_n718), .B2(new_n719), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n704), .B(new_n714), .C1(new_n717), .C2(new_n477), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(KEYINPUT112), .A3(new_n725), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n544), .B1(new_n733), .B2(new_n473), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n586), .A2(new_n702), .A3(new_n722), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n473), .A3(new_n544), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1328gat));
  OAI21_X1  g540(.A(G36gat), .B1(new_n733), .B2(new_n413), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n735), .A2(G36gat), .A3(new_n413), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT114), .B(KEYINPUT46), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(G1329gat));
  NOR3_X1   g545(.A1(new_n735), .A2(new_n691), .A3(new_n540), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n721), .A2(new_n484), .A3(new_n726), .ZN(new_n750));
  INV_X1    g549(.A(new_n540), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n484), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n727), .A2(new_n732), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n747), .B1(new_n754), .B2(new_n540), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g555(.A1(new_n735), .A2(G50gat), .A3(new_n269), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n721), .A2(new_n269), .A3(new_n726), .ZN(new_n760));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n727), .A2(new_n732), .A3(new_n522), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n763), .A2(KEYINPUT115), .A3(G50gat), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT115), .B1(new_n763), .B2(G50gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n757), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n766), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g566(.A(new_n724), .ZN(new_n768));
  INV_X1    g567(.A(new_n657), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n702), .A2(new_n768), .A3(new_n769), .A4(new_n677), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n718), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n473), .B(KEYINPUT116), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(new_n640), .Z(G1332gat));
  NOR2_X1   g573(.A1(new_n771), .A2(new_n413), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  AND2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n775), .B2(new_n776), .ZN(G1333gat));
  NOR3_X1   g578(.A1(new_n771), .A2(G71gat), .A3(new_n691), .ZN(new_n780));
  INV_X1    g579(.A(new_n771), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n753), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(G71gat), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n522), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g585(.A1(new_n718), .A2(new_n724), .A3(new_n769), .A4(new_n702), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT51), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n677), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n591), .A3(new_n682), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n676), .A2(new_n724), .A3(new_n769), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n721), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n473), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1336gat));
  AOI21_X1  g594(.A(new_n590), .B1(new_n792), .B2(new_n412), .ZN(new_n796));
  INV_X1    g595(.A(new_n788), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n677), .A2(G92gat), .A3(new_n413), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT117), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n801), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n800), .A2(new_n801), .B1(new_n796), .B2(new_n803), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n793), .B2(new_n484), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n677), .A2(G99gat), .A3(new_n691), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n269), .A2(G106gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT118), .B1(new_n789), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n793), .B2(new_n269), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g612(.A1(new_n575), .A2(new_n576), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n529), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n676), .A2(new_n580), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n663), .A2(new_n662), .A3(new_n666), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n818), .A2(new_n667), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n660), .B1(new_n667), .B2(new_n819), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT54), .B(new_n662), .C1(new_n663), .C2(new_n666), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT119), .B1(new_n824), .B2(new_n660), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n820), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n675), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  AOI211_X1 g627(.A(new_n828), .B(new_n820), .C1(new_n823), .C2(new_n825), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n768), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n702), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n580), .A3(new_n816), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n629), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n769), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n678), .A2(new_n768), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n772), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n413), .A3(new_n377), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n768), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n835), .A2(new_n837), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n473), .A2(new_n412), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n842), .A2(new_n522), .A3(new_n691), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n585), .A2(new_n325), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n840), .B2(new_n676), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n842), .A2(new_n522), .A3(new_n844), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n677), .A2(new_n323), .A3(new_n691), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n318), .A2(new_n319), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n845), .A2(new_n853), .A3(new_n657), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n840), .B2(new_n657), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1342gat));
  NOR3_X1   g657(.A1(new_n839), .A2(G134gat), .A3(new_n629), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n702), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G134gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n753), .A2(new_n844), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n835), .A2(new_n837), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n522), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n830), .A2(new_n584), .A3(new_n581), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n869), .A2(new_n817), .B1(new_n628), .B2(new_n623), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n769), .B1(new_n834), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n836), .B1(new_n871), .B2(KEYINPUT121), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n769), .C1(new_n834), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n269), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n865), .B1(new_n868), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n216), .B1(new_n879), .B2(new_n768), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n753), .A2(new_n412), .A3(new_n269), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n838), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n585), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n877), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n872), .B2(new_n874), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n864), .B1(new_n867), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n585), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT122), .B1(new_n882), .B2(new_n884), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n838), .A2(new_n892), .A3(new_n881), .A4(new_n883), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT123), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n890), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n702), .A2(new_n769), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n585), .A4(new_n677), .ZN(new_n900));
  INV_X1    g699(.A(new_n585), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT124), .B1(new_n678), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n871), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n522), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n904), .A2(new_n905), .B1(new_n842), .B2(new_n887), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT125), .B(KEYINPUT57), .C1(new_n903), .C2(new_n522), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n864), .A2(new_n676), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT59), .B(G148gat), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n882), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n214), .A3(new_n676), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n214), .B1(new_n879), .B2(new_n676), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n910), .B(new_n912), .C1(KEYINPUT59), .C2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n889), .B2(new_n769), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n769), .A2(G155gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n882), .B2(new_n916), .ZN(G1346gat));
  AOI21_X1  g716(.A(G162gat), .B1(new_n911), .B2(new_n702), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n702), .A2(G162gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n879), .B2(new_n919), .ZN(G1347gat));
  NAND2_X1  g719(.A1(new_n772), .A2(new_n412), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n691), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n866), .A2(new_n269), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n309), .A3(new_n585), .ZN(new_n924));
  NOR4_X1   g723(.A1(new_n842), .A2(new_n682), .A3(new_n413), .A4(new_n376), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n768), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n926), .B2(new_n309), .ZN(G1348gat));
  NOR3_X1   g726(.A1(new_n923), .A2(new_n310), .A3(new_n677), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n676), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n310), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n274), .A2(G183gat), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n925), .A2(new_n931), .A3(new_n276), .A4(new_n657), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n281), .A2(G183gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n923), .A2(new_n769), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n923), .B2(new_n629), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n925), .A2(new_n302), .A3(new_n702), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n921), .A2(new_n753), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n585), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n942), .B(new_n944), .C1(new_n906), .C2(new_n907), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n753), .A2(new_n413), .A3(new_n269), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n866), .A2(new_n473), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(new_n724), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(KEYINPUT126), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1352gat));
  OR2_X1    g752(.A1(new_n906), .A2(new_n907), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n676), .A3(new_n942), .ZN(new_n955));
  XOR2_X1   g754(.A(KEYINPUT127), .B(G204gat), .Z(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n947), .A2(new_n677), .A3(new_n956), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  OR3_X1    g759(.A1(new_n947), .A2(G211gat), .A3(new_n769), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n657), .B(new_n942), .C1(new_n906), .C2(new_n907), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NAND3_X1  g764(.A1(new_n954), .A2(new_n702), .A3(new_n942), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G218gat), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n947), .A2(G218gat), .A3(new_n629), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1355gat));
endmodule


