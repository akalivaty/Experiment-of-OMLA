

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  NOR2_X1 U321 ( .A1(n531), .A2(n469), .ZN(n558) );
  XNOR2_X1 U322 ( .A(n303), .B(n302), .ZN(n518) );
  XOR2_X1 U323 ( .A(n419), .B(n418), .Z(n289) );
  XOR2_X1 U324 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n290) );
  XNOR2_X1 U325 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n292) );
  XNOR2_X1 U326 ( .A(n387), .B(n292), .ZN(n295) );
  XNOR2_X1 U327 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U329 ( .A1(n578), .A2(n408), .ZN(n409) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n471) );
  XNOR2_X1 U331 ( .A(KEYINPUT38), .B(n446), .ZN(n499) );
  XNOR2_X1 U332 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U333 ( .A(n447), .B(G36GAT), .ZN(n448) );
  XNOR2_X1 U334 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(n449), .B(n448), .ZN(G1329GAT) );
  XOR2_X1 U336 ( .A(G183GAT), .B(KEYINPUT86), .Z(n327) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n290), .B(n291), .ZN(n387) );
  XOR2_X1 U339 ( .A(G169GAT), .B(G8GAT), .Z(n431) );
  XNOR2_X1 U340 ( .A(G36GAT), .B(n431), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(G204GAT), .ZN(n294) );
  XOR2_X1 U342 ( .A(n295), .B(n294), .Z(n300) );
  XOR2_X1 U343 ( .A(G211GAT), .B(KEYINPUT21), .Z(n297) );
  XNOR2_X1 U344 ( .A(G197GAT), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n378) );
  XNOR2_X1 U346 ( .A(G176GAT), .B(G92GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n298), .B(G64GAT), .ZN(n411) );
  XNOR2_X1 U348 ( .A(n378), .B(n411), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n327), .B(n301), .Z(n303) );
  NAND2_X1 U351 ( .A1(G226GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT73), .Z(n305) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G36GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n443) );
  INV_X1 U357 ( .A(n443), .ZN(n311) );
  XOR2_X1 U358 ( .A(KEYINPUT67), .B(KEYINPUT84), .Z(n309) );
  XNOR2_X1 U359 ( .A(G162GAT), .B(KEYINPUT85), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n324) );
  XOR2_X1 U362 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n313) );
  XNOR2_X1 U363 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U365 ( .A(KEYINPUT11), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .Z(n414) );
  XOR2_X1 U370 ( .A(n414), .B(G106GAT), .Z(n319) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(G134GAT), .B(n320), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n470) );
  XNOR2_X1 U376 ( .A(n470), .B(KEYINPUT36), .ZN(n578) );
  XOR2_X1 U377 ( .A(G78GAT), .B(G211GAT), .Z(n326) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(G71GAT), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U380 ( .A(n328), .B(n327), .Z(n330) );
  XNOR2_X1 U381 ( .A(G22GAT), .B(G155GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U383 ( .A(KEYINPUT88), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U386 ( .A(n334), .B(n333), .Z(n338) );
  XNOR2_X1 U387 ( .A(G15GAT), .B(G1GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n335), .B(KEYINPUT74), .ZN(n437) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(KEYINPUT77), .ZN(n410) );
  XNOR2_X1 U391 ( .A(n437), .B(n410), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n340) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT87), .B(n341), .Z(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n575) );
  INV_X1 U398 ( .A(n575), .ZN(n475) );
  XOR2_X1 U399 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n345) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n364) );
  XOR2_X1 U402 ( .A(G127GAT), .B(KEYINPUT0), .Z(n347) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(G134GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n385) );
  XOR2_X1 U405 ( .A(G155GAT), .B(KEYINPUT2), .Z(n349) );
  XNOR2_X1 U406 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n365) );
  XNOR2_X1 U408 ( .A(n385), .B(n365), .ZN(n362) );
  XOR2_X1 U409 ( .A(G85GAT), .B(G120GAT), .Z(n351) );
  XNOR2_X1 U410 ( .A(G29GAT), .B(G141GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U412 ( .A(KEYINPUT6), .B(G57GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G148GAT), .B(KEYINPUT93), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n357) );
  NAND2_X1 U417 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U419 ( .A(KEYINPUT94), .B(n358), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n562) );
  XOR2_X1 U423 ( .A(KEYINPUT24), .B(n365), .Z(n367) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U426 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n369) );
  XNOR2_X1 U427 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U429 ( .A(n371), .B(n370), .Z(n376) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(G22GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n372), .B(G141GAT), .ZN(n438) );
  XOR2_X1 U432 ( .A(G78GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U433 ( .A(G106GAT), .B(G204GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n421) );
  XNOR2_X1 U435 ( .A(n438), .B(n421), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U437 ( .A(n378), .B(n377), .Z(n466) );
  XNOR2_X1 U438 ( .A(n466), .B(KEYINPUT28), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n379), .B(KEYINPUT68), .ZN(n530) );
  XOR2_X1 U440 ( .A(n518), .B(KEYINPUT99), .Z(n380) );
  XNOR2_X1 U441 ( .A(KEYINPUT27), .B(n380), .ZN(n526) );
  NOR2_X1 U442 ( .A1(n530), .A2(n526), .ZN(n395) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n382) );
  XNOR2_X1 U444 ( .A(G15GAT), .B(KEYINPUT89), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n394) );
  XOR2_X1 U446 ( .A(G183GAT), .B(G176GAT), .Z(n384) );
  NAND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n386) );
  XOR2_X1 U449 ( .A(n386), .B(n385), .Z(n389) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U452 ( .A(G120GAT), .B(G71GAT), .Z(n415) );
  XOR2_X1 U453 ( .A(n390), .B(n415), .Z(n392) );
  XNOR2_X1 U454 ( .A(G43GAT), .B(G99GAT), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n531) );
  NAND2_X1 U457 ( .A1(n395), .A2(n531), .ZN(n396) );
  NOR2_X1 U458 ( .A1(n562), .A2(n396), .ZN(n397) );
  XOR2_X1 U459 ( .A(n397), .B(KEYINPUT100), .Z(n407) );
  NOR2_X1 U460 ( .A1(n518), .A2(n531), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n398), .B(KEYINPUT102), .ZN(n399) );
  NOR2_X1 U462 ( .A1(n466), .A2(n399), .ZN(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT25), .B(n400), .ZN(n404) );
  NAND2_X1 U464 ( .A1(n531), .A2(n466), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n401), .B(KEYINPUT26), .ZN(n565) );
  NOR2_X1 U466 ( .A1(n565), .A2(n526), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT101), .ZN(n403) );
  NAND2_X1 U468 ( .A1(n404), .A2(n403), .ZN(n405) );
  NAND2_X1 U469 ( .A1(n562), .A2(n405), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n407), .A2(n406), .ZN(n477) );
  NAND2_X1 U471 ( .A1(n475), .A2(n477), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT37), .B(n409), .Z(n516) );
  XOR2_X1 U473 ( .A(n411), .B(n410), .Z(n427) );
  XOR2_X1 U474 ( .A(KEYINPUT78), .B(KEYINPUT81), .Z(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT82), .B(KEYINPUT80), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U477 ( .A(KEYINPUT79), .B(KEYINPUT32), .Z(n417) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  NAND2_X1 U480 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n289), .B(n420), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n421), .B(KEYINPUT31), .ZN(n423) );
  INV_X1 U483 ( .A(KEYINPUT33), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n570) );
  XOR2_X1 U485 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n430), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(n431), .B(G113GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n442) );
  XOR2_X1 U491 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n435) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(KEYINPUT75), .Z(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n501) );
  INV_X1 U499 ( .A(n501), .ZN(n566) );
  XNOR2_X1 U500 ( .A(KEYINPUT76), .B(n566), .ZN(n551) );
  NAND2_X1 U501 ( .A1(n570), .A2(n551), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT83), .ZN(n480) );
  NAND2_X1 U503 ( .A1(n516), .A2(n480), .ZN(n446) );
  NOR2_X1 U504 ( .A1(n518), .A2(n499), .ZN(n449) );
  XNOR2_X1 U505 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT47), .B(KEYINPUT119), .Z(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT118), .B(KEYINPUT46), .ZN(n452) );
  XOR2_X1 U508 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n450) );
  XOR2_X1 U509 ( .A(n570), .B(n450), .Z(n543) );
  NAND2_X1 U510 ( .A1(n566), .A2(n543), .ZN(n451) );
  XOR2_X1 U511 ( .A(n452), .B(n451), .Z(n453) );
  NOR2_X1 U512 ( .A1(n575), .A2(n453), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n454), .A2(n470), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n475), .A2(n578), .ZN(n458) );
  XNOR2_X1 U516 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n459), .A2(n570), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n551), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT120), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT48), .B(n464), .ZN(n527) );
  NOR2_X1 U523 ( .A1(n518), .A2(n527), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT54), .ZN(n563) );
  INV_X1 U525 ( .A(n562), .ZN(n529) );
  NOR2_X1 U526 ( .A1(n529), .A2(n466), .ZN(n467) );
  AND2_X1 U527 ( .A1(n563), .A2(n467), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT55), .ZN(n469) );
  INV_X1 U529 ( .A(n470), .ZN(n549) );
  NAND2_X1 U530 ( .A1(n558), .A2(n549), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n472) );
  NOR2_X1 U532 ( .A1(n475), .A2(n549), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT16), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n502) );
  INV_X1 U535 ( .A(n502), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n490) );
  NOR2_X1 U537 ( .A1(n562), .A2(n490), .ZN(n482) );
  XNOR2_X1 U538 ( .A(KEYINPUT103), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n518), .A2(n490), .ZN(n485) );
  XNOR2_X1 U542 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U545 ( .A1(n531), .A2(n490), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT106), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  INV_X1 U549 ( .A(n530), .ZN(n522) );
  NOR2_X1 U550 ( .A1(n522), .A2(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT107), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U553 ( .A1(n499), .A2(n562), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT39), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n499), .A2(n531), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n522), .ZN(n500) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  XNOR2_X1 U563 ( .A(KEYINPUT112), .B(n543), .ZN(n553) );
  NAND2_X1 U564 ( .A1(n501), .A2(n553), .ZN(n514) );
  NOR2_X1 U565 ( .A1(n514), .A2(n502), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT113), .B(n503), .ZN(n511) );
  NOR2_X1 U567 ( .A1(n562), .A2(n511), .ZN(n504) );
  XOR2_X1 U568 ( .A(n504), .B(KEYINPUT42), .Z(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n518), .A2(n511), .ZN(n506) );
  XOR2_X1 U571 ( .A(KEYINPUT114), .B(n506), .Z(n507) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n531), .A2(n511), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n522), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  INV_X1 U580 ( .A(n514), .ZN(n515) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n521) );
  NOR2_X1 U582 ( .A1(n562), .A2(n521), .ZN(n517) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n521), .ZN(n519) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n521), .ZN(n520) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n520), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT117), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n541) );
  OR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n541), .A2(n532), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n538), .A2(n551), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n538), .A2(n553), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n575), .A2(n538), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n549), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n565), .A2(n541), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n548), .A2(n566), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U611 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n575), .A2(n548), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT121), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n558), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n575), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n572) );
  INV_X1 U636 ( .A(n574), .ZN(n577) );
  OR2_X1 U637 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

