

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834;

  BUF_X1 U374 ( .A(n833), .Z(n351) );
  BUF_X1 U375 ( .A(n798), .Z(n352) );
  OR2_X1 U376 ( .A1(n799), .A2(n629), .ZN(n437) );
  XNOR2_X1 U377 ( .A(n466), .B(n390), .ZN(n798) );
  XNOR2_X1 U378 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U379 ( .A(KEYINPUT110), .ZN(n354) );
  BUF_X1 U380 ( .A(n686), .Z(n432) );
  XNOR2_X1 U381 ( .A(n571), .B(n570), .ZN(n610) );
  OR2_X1 U382 ( .A1(n721), .A2(n699), .ZN(n571) );
  NAND2_X1 U383 ( .A1(n735), .A2(G475), .ZN(n729) );
  AND2_X2 U384 ( .A1(n706), .A2(n365), .ZN(n735) );
  NAND2_X1 U385 ( .A1(n735), .A2(G472), .ZN(n710) );
  NAND2_X2 U386 ( .A1(n395), .A2(n468), .ZN(n690) );
  NAND2_X2 U387 ( .A1(n442), .A2(n443), .ZN(n732) );
  XNOR2_X2 U388 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X2 U389 ( .A(n627), .B(n438), .ZN(n785) );
  NAND2_X1 U390 ( .A1(n735), .A2(G210), .ZN(n723) );
  XNOR2_X2 U391 ( .A(n727), .B(n726), .ZN(n728) );
  AND2_X2 U392 ( .A1(n456), .A2(n451), .ZN(n441) );
  NAND2_X1 U393 ( .A1(n353), .A2(n357), .ZN(n356) );
  INV_X1 U394 ( .A(n798), .ZN(n353) );
  OR2_X1 U395 ( .A1(n768), .A2(n771), .ZN(n355) );
  NAND2_X2 U396 ( .A1(n364), .A2(n467), .ZN(n363) );
  XNOR2_X2 U397 ( .A(n685), .B(KEYINPUT6), .ZN(n665) );
  XNOR2_X1 U398 ( .A(n356), .B(n391), .ZN(n400) );
  AND2_X2 U399 ( .A1(n403), .A2(n409), .ZN(n402) );
  XNOR2_X1 U400 ( .A(KEYINPUT81), .B(n506), .ZN(n573) );
  XOR2_X1 U401 ( .A(n690), .B(KEYINPUT100), .Z(n357) );
  XOR2_X1 U402 ( .A(n632), .B(n631), .Z(n359) );
  NOR2_X1 U403 ( .A1(n792), .A2(n352), .ZN(n360) );
  AND2_X2 U404 ( .A1(n376), .A2(n375), .ZN(n361) );
  NAND2_X2 U405 ( .A1(n405), .A2(n402), .ZN(n408) );
  NOR2_X2 U406 ( .A1(G953), .A2(G237), .ZN(n505) );
  INV_X1 U407 ( .A(KEYINPUT89), .ZN(n380) );
  NAND2_X1 U408 ( .A1(n682), .A2(n362), .ZN(n674) );
  XNOR2_X1 U409 ( .A(n435), .B(n633), .ZN(n718) );
  NAND2_X1 U410 ( .A1(n359), .A2(n433), .ZN(n435) );
  NOR2_X2 U411 ( .A1(n626), .A2(n601), .ZN(n759) );
  OR2_X1 U412 ( .A1(n727), .A2(G902), .ZN(n434) );
  OR2_X2 U413 ( .A1(n383), .A2(n454), .ZN(n453) );
  INV_X1 U414 ( .A(KEYINPUT42), .ZN(n436) );
  XNOR2_X1 U415 ( .A(n705), .B(n704), .ZN(n364) );
  NAND2_X1 U416 ( .A1(n368), .A2(n367), .ZN(n366) );
  AND2_X1 U417 ( .A1(n664), .A2(KEYINPUT44), .ZN(n673) );
  NAND2_X1 U418 ( .A1(n444), .A2(n445), .ZN(n442) );
  AND2_X1 U419 ( .A1(n446), .A2(n447), .ZN(n443) );
  INV_X1 U420 ( .A(n716), .ZN(n362) );
  OR2_X1 U421 ( .A1(n629), .A2(n388), .ZN(n620) );
  XNOR2_X1 U422 ( .A(n635), .B(n614), .ZN(n615) );
  INV_X1 U423 ( .A(n398), .ZN(n477) );
  AND2_X1 U424 ( .A1(n394), .A2(n470), .ZN(n396) );
  NAND2_X1 U425 ( .A1(n479), .A2(n478), .ZN(n398) );
  XNOR2_X1 U426 ( .A(n383), .B(n708), .ZN(n709) );
  XNOR2_X1 U427 ( .A(n434), .B(G475), .ZN(n586) );
  NOR2_X1 U428 ( .A1(G902), .A2(n739), .ZN(n597) );
  XNOR2_X1 U429 ( .A(n568), .B(n811), .ZN(n721) );
  XNOR2_X1 U430 ( .A(n533), .B(G902), .ZN(n699) );
  XNOR2_X1 U431 ( .A(G113), .B(G104), .ZN(n581) );
  XNOR2_X2 U432 ( .A(n363), .B(KEYINPUT82), .ZN(n706) );
  NAND2_X1 U433 ( .A1(n369), .A2(n366), .ZN(n365) );
  INV_X1 U434 ( .A(n385), .ZN(n367) );
  NAND2_X1 U435 ( .A1(n467), .A2(n492), .ZN(n368) );
  XNOR2_X2 U436 ( .A(n697), .B(KEYINPUT45), .ZN(n467) );
  NAND2_X1 U437 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U438 ( .A1(n490), .A2(n826), .ZN(n370) );
  NAND2_X1 U439 ( .A1(n491), .A2(n385), .ZN(n371) );
  XNOR2_X2 U440 ( .A(n372), .B(n634), .ZN(n703) );
  NAND2_X2 U441 ( .A1(n361), .A2(n373), .ZN(n372) );
  NOR2_X2 U442 ( .A1(n374), .A2(n422), .ZN(n373) );
  NAND2_X1 U443 ( .A1(n419), .A2(n417), .ZN(n374) );
  NAND2_X1 U444 ( .A1(n381), .A2(n425), .ZN(n375) );
  NAND2_X1 U445 ( .A1(n379), .A2(n426), .ZN(n376) );
  NAND2_X1 U446 ( .A1(n652), .A2(n651), .ZN(n482) );
  XNOR2_X2 U447 ( .A(n521), .B(n520), .ZN(n587) );
  XNOR2_X1 U448 ( .A(n377), .B(n378), .ZN(n686) );
  NOR2_X1 U449 ( .A1(n744), .A2(G902), .ZN(n377) );
  XOR2_X1 U450 ( .A(KEYINPUT73), .B(G469), .Z(n378) );
  NOR2_X1 U451 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U452 ( .A(n408), .B(n380), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n408), .B(KEYINPUT89), .ZN(n381) );
  NOR2_X1 U454 ( .A1(n718), .A2(KEYINPUT46), .ZN(n420) );
  AND2_X2 U455 ( .A1(n626), .A2(n601), .ZN(n761) );
  XNOR2_X1 U456 ( .A(n555), .B(KEYINPUT83), .ZN(n382) );
  XNOR2_X1 U457 ( .A(n555), .B(KEYINPUT83), .ZN(n630) );
  XNOR2_X1 U458 ( .A(n519), .B(n510), .ZN(n383) );
  XNOR2_X1 U459 ( .A(n519), .B(n510), .ZN(n707) );
  AND2_X1 U460 ( .A1(n646), .A2(n472), .ZN(n471) );
  NOR2_X1 U461 ( .A1(n628), .A2(KEYINPUT19), .ZN(n475) );
  AND2_X1 U462 ( .A1(n461), .A2(n389), .ZN(n460) );
  NAND2_X1 U463 ( .A1(n418), .A2(n426), .ZN(n417) );
  NAND2_X1 U464 ( .A1(n420), .A2(n421), .ZN(n419) );
  INV_X1 U465 ( .A(n624), .ZN(n418) );
  NAND2_X1 U466 ( .A1(n424), .A2(n423), .ZN(n422) );
  XNOR2_X1 U467 ( .A(KEYINPUT3), .B(G119), .ZN(n500) );
  NAND2_X1 U468 ( .A1(n495), .A2(n493), .ZN(n492) );
  NAND2_X1 U469 ( .A1(n699), .A2(n494), .ZN(n493) );
  NAND2_X1 U470 ( .A1(n496), .A2(KEYINPUT64), .ZN(n495) );
  NAND2_X1 U471 ( .A1(KEYINPUT2), .A2(KEYINPUT64), .ZN(n494) );
  NAND2_X1 U472 ( .A1(n785), .A2(n784), .ZN(n788) );
  INV_X1 U473 ( .A(G237), .ZN(n512) );
  INV_X1 U474 ( .A(G902), .ZN(n513) );
  NAND2_X1 U475 ( .A1(G472), .A2(n513), .ZN(n454) );
  NAND2_X1 U476 ( .A1(n511), .A2(G902), .ZN(n455) );
  INV_X1 U477 ( .A(KEYINPUT92), .ZN(n704) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n799) );
  INV_X1 U479 ( .A(KEYINPUT41), .ZN(n415) );
  NAND2_X1 U480 ( .A1(n785), .A2(n414), .ZN(n416) );
  NOR2_X1 U481 ( .A1(n787), .A2(n628), .ZN(n414) );
  NAND2_X1 U482 ( .A1(n473), .A2(n477), .ZN(n468) );
  AND2_X1 U483 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U484 ( .A1(n474), .A2(n649), .ZN(n473) );
  INV_X1 U485 ( .A(n767), .ZN(n413) );
  INV_X1 U486 ( .A(n685), .ZN(n774) );
  INV_X1 U487 ( .A(KEYINPUT71), .ZN(n426) );
  INV_X1 U488 ( .A(KEYINPUT15), .ZN(n533) );
  OR2_X1 U489 ( .A1(n771), .A2(n605), .ZN(n611) );
  NOR2_X1 U490 ( .A1(n628), .A2(n452), .ZN(n451) );
  INV_X1 U491 ( .A(KEYINPUT30), .ZN(n457) );
  XNOR2_X1 U492 ( .A(G113), .B(G137), .ZN(n504) );
  XNOR2_X1 U493 ( .A(KEYINPUT104), .B(KEYINPUT5), .ZN(n503) );
  XNOR2_X1 U494 ( .A(G131), .B(G134), .ZN(n820) );
  XNOR2_X1 U495 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n501) );
  XNOR2_X1 U496 ( .A(G116), .B(KEYINPUT74), .ZN(n499) );
  XNOR2_X1 U497 ( .A(G122), .B(G107), .ZN(n588) );
  XNOR2_X1 U498 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n563) );
  NAND2_X1 U499 ( .A1(G234), .A2(G237), .ZN(n540) );
  INV_X1 U500 ( .A(KEYINPUT38), .ZN(n438) );
  OR2_X1 U501 ( .A1(n646), .A2(n472), .ZN(n470) );
  NOR2_X1 U502 ( .A1(n627), .A2(n572), .ZN(n487) );
  NAND2_X1 U503 ( .A1(n628), .A2(KEYINPUT19), .ZN(n478) );
  XOR2_X1 U504 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n593) );
  XNOR2_X1 U505 ( .A(G116), .B(KEYINPUT108), .ZN(n592) );
  XOR2_X1 U506 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n579) );
  XNOR2_X1 U507 ( .A(KEYINPUT107), .B(KEYINPUT11), .ZN(n578) );
  XOR2_X1 U508 ( .A(KEYINPUT12), .B(G122), .Z(n575) );
  XNOR2_X1 U509 ( .A(n580), .B(n458), .ZN(n582) );
  XNOR2_X1 U510 ( .A(n581), .B(n459), .ZN(n458) );
  INV_X1 U511 ( .A(G140), .ZN(n459) );
  XNOR2_X1 U512 ( .A(G137), .B(G140), .ZN(n531) );
  XNOR2_X1 U513 ( .A(G110), .B(G104), .ZN(n514) );
  XNOR2_X1 U514 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n556) );
  NAND2_X1 U515 ( .A1(n358), .A2(n481), .ZN(n480) );
  INV_X1 U516 ( .A(n655), .ZN(n481) );
  NOR2_X1 U517 ( .A1(n658), .A2(n657), .ZN(n444) );
  AND2_X2 U518 ( .A1(n449), .A2(n428), .ZN(n685) );
  NOR2_X1 U519 ( .A1(n829), .A2(G952), .ZN(n747) );
  NOR2_X1 U520 ( .A1(n386), .A2(n427), .ZN(n803) );
  NAND2_X1 U521 ( .A1(n639), .A2(n439), .ZN(n715) );
  XNOR2_X1 U522 ( .A(n691), .B(KEYINPUT31), .ZN(n412) );
  BUF_X1 U523 ( .A(n759), .Z(n433) );
  OR2_X1 U524 ( .A1(n658), .A2(n655), .ZN(n684) );
  AND2_X1 U525 ( .A1(n476), .A2(n784), .ZN(n384) );
  AND2_X1 U526 ( .A1(n492), .A2(n392), .ZN(n385) );
  INV_X1 U527 ( .A(KEYINPUT64), .ZN(n700) );
  AND2_X1 U528 ( .A1(n497), .A2(n698), .ZN(n386) );
  AND2_X1 U529 ( .A1(n627), .A2(n572), .ZN(n387) );
  AND2_X1 U530 ( .A1(n474), .A2(n477), .ZN(n388) );
  AND2_X1 U531 ( .A1(n695), .A2(n696), .ZN(n389) );
  INV_X1 U532 ( .A(n668), .ZN(n488) );
  AND2_X1 U533 ( .A1(n599), .A2(n601), .ZN(n668) );
  XOR2_X1 U534 ( .A(KEYINPUT111), .B(KEYINPUT33), .Z(n390) );
  XOR2_X1 U535 ( .A(n667), .B(KEYINPUT78), .Z(n391) );
  AND2_X1 U536 ( .A1(n569), .A2(G214), .ZN(n628) );
  NAND2_X1 U537 ( .A1(n698), .A2(n700), .ZN(n392) );
  AND2_X1 U538 ( .A1(n699), .A2(KEYINPUT64), .ZN(n393) );
  NAND2_X1 U539 ( .A1(n476), .A2(n469), .ZN(n394) );
  NAND2_X1 U540 ( .A1(n398), .A2(n471), .ZN(n397) );
  XNOR2_X2 U541 ( .A(n399), .B(n670), .ZN(n719) );
  NAND2_X1 U542 ( .A1(n400), .A2(n668), .ZN(n399) );
  NAND2_X1 U543 ( .A1(n620), .A2(KEYINPUT47), .ZN(n409) );
  NAND2_X1 U544 ( .A1(n733), .A2(n404), .ZN(n403) );
  AND2_X1 U545 ( .A1(n603), .A2(n484), .ZN(n404) );
  NOR2_X1 U546 ( .A1(n603), .A2(n484), .ZN(n406) );
  NOR2_X1 U547 ( .A1(n733), .A2(n484), .ZN(n407) );
  NAND2_X1 U548 ( .A1(n411), .A2(n410), .ZN(n693) );
  INV_X1 U549 ( .A(n750), .ZN(n410) );
  INV_X1 U550 ( .A(n412), .ZN(n411) );
  NAND2_X1 U551 ( .A1(n412), .A2(n761), .ZN(n762) );
  NAND2_X1 U552 ( .A1(n412), .A2(n433), .ZN(n760) );
  NAND2_X1 U553 ( .A1(n685), .A2(n413), .ZN(n689) );
  INV_X1 U554 ( .A(n833), .ZN(n421) );
  NAND2_X1 U555 ( .A1(n718), .A2(KEYINPUT46), .ZN(n423) );
  NAND2_X1 U556 ( .A1(n833), .A2(KEYINPUT46), .ZN(n424) );
  AND2_X1 U557 ( .A1(n624), .A2(KEYINPUT71), .ZN(n425) );
  XNOR2_X2 U558 ( .A(n437), .B(n436), .ZN(n833) );
  INV_X1 U559 ( .A(n706), .ZN(n427) );
  BUF_X1 U560 ( .A(n735), .Z(n742) );
  NAND2_X1 U561 ( .A1(n441), .A2(n453), .ZN(n440) );
  BUF_X1 U562 ( .A(n456), .Z(n428) );
  XNOR2_X2 U563 ( .A(n429), .B(n600), .ZN(n733) );
  NAND2_X2 U564 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U565 ( .A1(n485), .A2(KEYINPUT112), .ZN(n430) );
  AND2_X2 U566 ( .A1(n489), .A2(n486), .ZN(n431) );
  XNOR2_X1 U567 ( .A(n440), .B(n457), .ZN(n554) );
  OR2_X2 U568 ( .A1(n665), .A2(n613), .ZN(n635) );
  INV_X1 U569 ( .A(n627), .ZN(n439) );
  XNOR2_X2 U570 ( .A(n562), .B(n498), .ZN(n519) );
  INV_X1 U571 ( .A(n480), .ZN(n445) );
  NAND2_X1 U572 ( .A1(n658), .A2(n657), .ZN(n446) );
  NAND2_X1 U573 ( .A1(n480), .A2(n657), .ZN(n447) );
  XNOR2_X2 U574 ( .A(n432), .B(KEYINPUT1), .ZN(n768) );
  INV_X1 U575 ( .A(n450), .ZN(n449) );
  NAND2_X1 U576 ( .A1(n453), .A2(n455), .ZN(n450) );
  INV_X1 U577 ( .A(n455), .ZN(n452) );
  NAND2_X1 U578 ( .A1(n707), .A2(n511), .ZN(n456) );
  XNOR2_X2 U579 ( .A(n539), .B(n538), .ZN(n771) );
  XNOR2_X2 U580 ( .A(n586), .B(KEYINPUT13), .ZN(n626) );
  NOR2_X2 U581 ( .A1(n759), .A2(n761), .ZN(n789) );
  INV_X1 U582 ( .A(n699), .ZN(n496) );
  XNOR2_X2 U583 ( .A(n549), .B(n548), .ZN(n770) );
  NAND2_X1 U584 ( .A1(n462), .A2(n460), .ZN(n697) );
  NAND2_X1 U585 ( .A1(n680), .A2(KEYINPUT93), .ZN(n461) );
  NAND2_X1 U586 ( .A1(n679), .A2(n463), .ZN(n462) );
  NAND2_X1 U587 ( .A1(n464), .A2(n678), .ZN(n463) );
  NAND2_X1 U588 ( .A1(n680), .A2(n675), .ZN(n464) );
  NOR2_X2 U589 ( .A1(n666), .A2(n768), .ZN(n466) );
  NAND2_X1 U590 ( .A1(n467), .A2(n393), .ZN(n490) );
  NAND2_X1 U591 ( .A1(n827), .A2(n467), .ZN(n497) );
  NAND2_X1 U592 ( .A1(n467), .A2(n829), .ZN(n810) );
  NAND2_X1 U593 ( .A1(n476), .A2(n475), .ZN(n474) );
  AND2_X1 U594 ( .A1(n471), .A2(n475), .ZN(n469) );
  INV_X1 U595 ( .A(n649), .ZN(n472) );
  INV_X1 U596 ( .A(n610), .ZN(n476) );
  NAND2_X1 U597 ( .A1(n610), .A2(KEYINPUT19), .ZN(n479) );
  XNOR2_X2 U598 ( .A(n482), .B(n654), .ZN(n658) );
  XNOR2_X2 U599 ( .A(n483), .B(G143), .ZN(n591) );
  XNOR2_X2 U600 ( .A(G128), .B(KEYINPUT87), .ZN(n483) );
  INV_X1 U601 ( .A(KEYINPUT88), .ZN(n484) );
  INV_X1 U602 ( .A(n382), .ZN(n485) );
  NOR2_X1 U603 ( .A1(n488), .A2(n487), .ZN(n486) );
  NAND2_X1 U604 ( .A1(n630), .A2(n387), .ZN(n489) );
  INV_X1 U605 ( .A(n826), .ZN(n491) );
  XNOR2_X2 U606 ( .A(n591), .B(KEYINPUT4), .ZN(n818) );
  XNOR2_X2 U607 ( .A(n818), .B(G101), .ZN(n562) );
  XNOR2_X1 U608 ( .A(n820), .B(G146), .ZN(n498) );
  XNOR2_X1 U609 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n502), .B(n501), .ZN(n566) );
  XNOR2_X1 U611 ( .A(n504), .B(n503), .ZN(n508) );
  INV_X1 U612 ( .A(n505), .ZN(n506) );
  NAND2_X1 U613 ( .A1(n573), .A2(G210), .ZN(n507) );
  XNOR2_X1 U614 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U615 ( .A(n566), .B(n509), .ZN(n510) );
  INV_X1 U616 ( .A(G472), .ZN(n511) );
  NAND2_X1 U617 ( .A1(n513), .A2(n512), .ZN(n569) );
  XNOR2_X1 U618 ( .A(n531), .B(n514), .ZN(n517) );
  INV_X4 U619 ( .A(G953), .ZN(n829) );
  NAND2_X1 U620 ( .A1(G227), .A2(n829), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n515), .B(G107), .ZN(n516) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U623 ( .A(n519), .B(n518), .ZN(n744) );
  XNOR2_X1 U624 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n521) );
  NAND2_X1 U625 ( .A1(n829), .A2(G234), .ZN(n520) );
  NAND2_X1 U626 ( .A1(n587), .A2(G221), .ZN(n529) );
  XNOR2_X1 U627 ( .A(G128), .B(G110), .ZN(n523) );
  XNOR2_X1 U628 ( .A(G119), .B(KEYINPUT101), .ZN(n522) );
  XNOR2_X1 U629 ( .A(n523), .B(n522), .ZN(n527) );
  XNOR2_X1 U630 ( .A(KEYINPUT24), .B(KEYINPUT77), .ZN(n525) );
  XNOR2_X1 U631 ( .A(KEYINPUT102), .B(KEYINPUT23), .ZN(n524) );
  XNOR2_X1 U632 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n532) );
  XNOR2_X1 U635 ( .A(G146), .B(G125), .ZN(n557) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n557), .B(n530), .ZN(n576) );
  XNOR2_X1 U638 ( .A(n576), .B(n531), .ZN(n822) );
  XNOR2_X1 U639 ( .A(n532), .B(n822), .ZN(n736) );
  OR2_X1 U640 ( .A1(n736), .A2(G902), .ZN(n539) );
  NAND2_X1 U641 ( .A1(n496), .A2(G234), .ZN(n534) );
  XNOR2_X1 U642 ( .A(n534), .B(KEYINPUT20), .ZN(n545) );
  NAND2_X1 U643 ( .A1(n545), .A2(G217), .ZN(n537) );
  XNOR2_X1 U644 ( .A(KEYINPUT84), .B(KEYINPUT103), .ZN(n535) );
  XNOR2_X1 U645 ( .A(n535), .B(KEYINPUT25), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(KEYINPUT97), .Z(n541) );
  XNOR2_X1 U648 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U649 ( .A1(G952), .A2(n542), .ZN(n796) );
  NOR2_X1 U650 ( .A1(G953), .A2(n796), .ZN(n643) );
  AND2_X1 U651 ( .A1(G902), .A2(n542), .ZN(n641) );
  NAND2_X1 U652 ( .A1(G953), .A2(n641), .ZN(n543) );
  NOR2_X1 U653 ( .A1(n543), .A2(G900), .ZN(n544) );
  OR2_X1 U654 ( .A1(n643), .A2(n544), .ZN(n550) );
  INV_X1 U655 ( .A(n545), .ZN(n547) );
  INV_X1 U656 ( .A(G221), .ZN(n546) );
  OR2_X1 U657 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U658 ( .A(KEYINPUT21), .ZN(n548) );
  NAND2_X1 U659 ( .A1(n550), .A2(n770), .ZN(n604) );
  INV_X1 U660 ( .A(n604), .ZN(n551) );
  NAND2_X1 U661 ( .A1(n771), .A2(n551), .ZN(n552) );
  NOR2_X1 U662 ( .A1(n686), .A2(n552), .ZN(n553) );
  NAND2_X1 U663 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n557), .B(n556), .ZN(n560) );
  NAND2_X1 U665 ( .A1(n829), .A2(G224), .ZN(n558) );
  XNOR2_X1 U666 ( .A(n558), .B(KEYINPUT96), .ZN(n559) );
  XNOR2_X1 U667 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U668 ( .A(n562), .B(n561), .ZN(n568) );
  XNOR2_X1 U669 ( .A(n581), .B(n588), .ZN(n565) );
  XNOR2_X1 U670 ( .A(n563), .B(G110), .ZN(n564) );
  XNOR2_X1 U671 ( .A(n565), .B(n564), .ZN(n567) );
  XNOR2_X1 U672 ( .A(n567), .B(n566), .ZN(n811) );
  NAND2_X1 U673 ( .A1(n569), .A2(G210), .ZN(n570) );
  INV_X1 U674 ( .A(n610), .ZN(n627) );
  INV_X1 U675 ( .A(KEYINPUT112), .ZN(n572) );
  NAND2_X1 U676 ( .A1(n573), .A2(G214), .ZN(n574) );
  XNOR2_X1 U677 ( .A(n575), .B(n574), .ZN(n577) );
  XNOR2_X1 U678 ( .A(n577), .B(n576), .ZN(n585) );
  XNOR2_X1 U679 ( .A(n579), .B(n578), .ZN(n583) );
  XNOR2_X1 U680 ( .A(G143), .B(G131), .ZN(n580) );
  XNOR2_X1 U681 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U682 ( .A(n585), .B(n584), .ZN(n727) );
  INV_X1 U683 ( .A(n626), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n587), .A2(G217), .ZN(n590) );
  XNOR2_X1 U685 ( .A(n588), .B(G134), .ZN(n589) );
  XNOR2_X1 U686 ( .A(n590), .B(n589), .ZN(n596) );
  XNOR2_X1 U687 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U688 ( .A(n591), .B(n594), .ZN(n595) );
  XNOR2_X1 U689 ( .A(n596), .B(n595), .ZN(n739) );
  XOR2_X1 U690 ( .A(n597), .B(KEYINPUT109), .Z(n598) );
  XNOR2_X1 U691 ( .A(n598), .B(G478), .ZN(n625) );
  INV_X1 U692 ( .A(n625), .ZN(n601) );
  INV_X1 U693 ( .A(KEYINPUT113), .ZN(n600) );
  NAND2_X1 U694 ( .A1(n789), .A2(KEYINPUT47), .ZN(n602) );
  XNOR2_X1 U695 ( .A(n602), .B(KEYINPUT90), .ZN(n603) );
  XNOR2_X1 U696 ( .A(n604), .B(KEYINPUT72), .ZN(n605) );
  OR2_X1 U697 ( .A1(n774), .A2(n611), .ZN(n607) );
  INV_X1 U698 ( .A(KEYINPUT28), .ZN(n606) );
  XNOR2_X1 U699 ( .A(n607), .B(n606), .ZN(n609) );
  INV_X1 U700 ( .A(n432), .ZN(n608) );
  NAND2_X1 U701 ( .A1(n609), .A2(n608), .ZN(n629) );
  INV_X1 U702 ( .A(n611), .ZN(n612) );
  NAND2_X1 U703 ( .A1(n759), .A2(n612), .ZN(n613) );
  INV_X1 U704 ( .A(KEYINPUT114), .ZN(n614) );
  NAND2_X1 U705 ( .A1(n615), .A2(n384), .ZN(n617) );
  INV_X1 U706 ( .A(KEYINPUT36), .ZN(n616) );
  XNOR2_X1 U707 ( .A(n617), .B(n616), .ZN(n619) );
  INV_X1 U708 ( .A(n768), .ZN(n618) );
  NAND2_X1 U709 ( .A1(n619), .A2(n618), .ZN(n764) );
  INV_X1 U710 ( .A(n620), .ZN(n757) );
  XNOR2_X1 U711 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n621) );
  NOR2_X1 U712 ( .A1(n789), .A2(n621), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n757), .A2(n622), .ZN(n623) );
  AND2_X1 U714 ( .A1(n764), .A2(n623), .ZN(n624) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n787) );
  INV_X1 U716 ( .A(n628), .ZN(n784) );
  NAND2_X1 U717 ( .A1(n382), .A2(n785), .ZN(n632) );
  INV_X1 U718 ( .A(KEYINPUT39), .ZN(n631) );
  INV_X1 U719 ( .A(KEYINPUT40), .ZN(n633) );
  INV_X1 U720 ( .A(KEYINPUT48), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n359), .A2(n761), .ZN(n714) );
  INV_X1 U722 ( .A(n635), .ZN(n637) );
  AND2_X1 U723 ( .A1(n768), .A2(n784), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT43), .ZN(n639) );
  AND2_X1 U726 ( .A1(n714), .A2(n715), .ZN(n701) );
  NAND2_X1 U727 ( .A1(n703), .A2(n701), .ZN(n640) );
  XNOR2_X2 U728 ( .A(n640), .B(KEYINPUT91), .ZN(n826) );
  NOR2_X1 U729 ( .A1(G898), .A2(n829), .ZN(n812) );
  NAND2_X1 U730 ( .A1(n812), .A2(n641), .ZN(n642) );
  XOR2_X1 U731 ( .A(KEYINPUT98), .B(n642), .Z(n644) );
  NOR2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U733 ( .A(n645), .B(KEYINPUT99), .ZN(n646) );
  XNOR2_X1 U734 ( .A(KEYINPUT94), .B(KEYINPUT0), .ZN(n648) );
  INV_X1 U735 ( .A(KEYINPUT67), .ZN(n647) );
  XNOR2_X1 U736 ( .A(n648), .B(n647), .ZN(n649) );
  INV_X1 U737 ( .A(n690), .ZN(n652) );
  INV_X1 U738 ( .A(n770), .ZN(n650) );
  NOR2_X1 U739 ( .A1(n787), .A2(n650), .ZN(n651) );
  INV_X1 U740 ( .A(KEYINPUT79), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n653), .B(KEYINPUT22), .ZN(n654) );
  INV_X1 U742 ( .A(n665), .ZN(n655) );
  INV_X1 U743 ( .A(KEYINPUT66), .ZN(n656) );
  XNOR2_X1 U744 ( .A(n656), .B(KEYINPUT32), .ZN(n657) );
  INV_X1 U745 ( .A(n658), .ZN(n662) );
  INV_X1 U746 ( .A(n771), .ZN(n659) );
  AND2_X1 U747 ( .A1(n774), .A2(n659), .ZN(n660) );
  AND2_X1 U748 ( .A1(n768), .A2(n660), .ZN(n661) );
  AND2_X1 U749 ( .A1(n662), .A2(n661), .ZN(n716) );
  INV_X1 U750 ( .A(KEYINPUT65), .ZN(n663) );
  NAND2_X1 U751 ( .A1(n674), .A2(n663), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n771), .A2(n770), .ZN(n767) );
  OR2_X2 U753 ( .A1(n665), .A2(n767), .ZN(n666) );
  XNOR2_X1 U754 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n667) );
  INV_X1 U755 ( .A(KEYINPUT85), .ZN(n669) );
  XNOR2_X1 U756 ( .A(n669), .B(KEYINPUT35), .ZN(n670) );
  INV_X1 U757 ( .A(KEYINPUT93), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n719), .A2(n671), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n679) );
  INV_X1 U760 ( .A(n674), .ZN(n675) );
  INV_X1 U761 ( .A(n719), .ZN(n680) );
  NOR2_X1 U762 ( .A1(KEYINPUT93), .A2(KEYINPUT65), .ZN(n677) );
  INV_X1 U763 ( .A(KEYINPUT44), .ZN(n676) );
  AND2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n678) );
  INV_X1 U765 ( .A(n732), .ZN(n682) );
  AND2_X1 U766 ( .A1(n362), .A2(KEYINPUT65), .ZN(n681) );
  NAND2_X1 U767 ( .A1(n682), .A2(n681), .ZN(n696) );
  NAND2_X1 U768 ( .A1(n768), .A2(n771), .ZN(n683) );
  OR2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n717) );
  OR2_X1 U770 ( .A1(n685), .A2(n767), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n687), .A2(n432), .ZN(n688) );
  AND2_X1 U772 ( .A1(n357), .A2(n688), .ZN(n750) );
  OR2_X1 U773 ( .A1(n768), .A2(n689), .ZN(n778) );
  OR2_X1 U774 ( .A1(n690), .A2(n778), .ZN(n691) );
  INV_X1 U775 ( .A(n789), .ZN(n692) );
  NAND2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U777 ( .A1(n717), .A2(n694), .ZN(n695) );
  INV_X1 U778 ( .A(KEYINPUT2), .ZN(n698) );
  AND2_X1 U779 ( .A1(n701), .A2(KEYINPUT2), .ZN(n702) );
  NAND2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n705) );
  XOR2_X1 U781 ( .A(KEYINPUT95), .B(KEYINPUT62), .Z(n708) );
  XNOR2_X1 U782 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X2 U783 ( .A1(n711), .A2(n747), .ZN(n713) );
  INV_X1 U784 ( .A(KEYINPUT63), .ZN(n712) );
  XNOR2_X1 U785 ( .A(n713), .B(n712), .ZN(G57) );
  XNOR2_X1 U786 ( .A(n714), .B(G134), .ZN(G36) );
  XNOR2_X1 U787 ( .A(n715), .B(G140), .ZN(G42) );
  XOR2_X1 U788 ( .A(G110), .B(n716), .Z(G12) );
  XNOR2_X1 U789 ( .A(n717), .B(G101), .ZN(G3) );
  XOR2_X1 U790 ( .A(G131), .B(n718), .Z(G33) );
  XOR2_X1 U791 ( .A(n719), .B(G122), .Z(G24) );
  XOR2_X1 U792 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n720) );
  XNOR2_X1 U793 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X2 U794 ( .A1(n724), .A2(n747), .ZN(n725) );
  XNOR2_X1 U795 ( .A(n725), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U796 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n726) );
  XNOR2_X1 U797 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X2 U798 ( .A1(n730), .A2(n747), .ZN(n731) );
  XNOR2_X1 U799 ( .A(n731), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U800 ( .A(n732), .B(G119), .Z(G21) );
  BUF_X1 U801 ( .A(n733), .Z(n734) );
  XNOR2_X1 U802 ( .A(n734), .B(G143), .ZN(G45) );
  NAND2_X1 U803 ( .A1(n742), .A2(G217), .ZN(n737) );
  XNOR2_X1 U804 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U805 ( .A1(n738), .A2(n747), .ZN(G66) );
  NAND2_X1 U806 ( .A1(n742), .A2(G478), .ZN(n740) );
  XNOR2_X1 U807 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U808 ( .A1(n741), .A2(n747), .ZN(G63) );
  NAND2_X1 U809 ( .A1(n742), .A2(G469), .ZN(n746) );
  XOR2_X1 U810 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n743) );
  XNOR2_X1 U811 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U812 ( .A(n746), .B(n745), .ZN(n748) );
  NOR2_X1 U813 ( .A1(n748), .A2(n747), .ZN(G54) );
  NAND2_X1 U814 ( .A1(n750), .A2(n433), .ZN(n749) );
  XNOR2_X1 U815 ( .A(n749), .B(G104), .ZN(G6) );
  XOR2_X1 U816 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n752) );
  NAND2_X1 U817 ( .A1(n750), .A2(n761), .ZN(n751) );
  XNOR2_X1 U818 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U819 ( .A(G107), .B(n753), .ZN(G9) );
  XOR2_X1 U820 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n755) );
  NAND2_X1 U821 ( .A1(n757), .A2(n761), .ZN(n754) );
  XNOR2_X1 U822 ( .A(n755), .B(n754), .ZN(n756) );
  XOR2_X1 U823 ( .A(G128), .B(n756), .Z(G30) );
  NAND2_X1 U824 ( .A1(n757), .A2(n433), .ZN(n758) );
  XNOR2_X1 U825 ( .A(n758), .B(G146), .ZN(G48) );
  XNOR2_X1 U826 ( .A(n760), .B(G113), .ZN(G15) );
  XNOR2_X1 U827 ( .A(n762), .B(KEYINPUT116), .ZN(n763) );
  XNOR2_X1 U828 ( .A(G116), .B(n763), .ZN(G18) );
  XOR2_X1 U829 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n766) );
  XOR2_X1 U830 ( .A(G125), .B(n764), .Z(n765) );
  XNOR2_X1 U831 ( .A(n766), .B(n765), .ZN(G27) );
  XOR2_X1 U832 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n806) );
  NAND2_X1 U833 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U834 ( .A(n769), .B(KEYINPUT50), .ZN(n777) );
  NOR2_X1 U835 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U836 ( .A(n772), .B(KEYINPUT49), .ZN(n773) );
  NAND2_X1 U837 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U838 ( .A(KEYINPUT118), .B(n775), .Z(n776) );
  NAND2_X1 U839 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U840 ( .A1(n779), .A2(n778), .ZN(n781) );
  XOR2_X1 U841 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n780) );
  XNOR2_X1 U842 ( .A(n781), .B(n780), .ZN(n782) );
  NOR2_X1 U843 ( .A1(n782), .A2(n799), .ZN(n783) );
  XNOR2_X1 U844 ( .A(n783), .B(KEYINPUT120), .ZN(n793) );
  NOR2_X1 U845 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U846 ( .A1(n787), .A2(n786), .ZN(n791) );
  NOR2_X1 U847 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U848 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U849 ( .A1(n793), .A2(n360), .ZN(n794) );
  XNOR2_X1 U850 ( .A(n794), .B(KEYINPUT52), .ZN(n795) );
  NOR2_X1 U851 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U852 ( .A(n797), .B(KEYINPUT121), .ZN(n801) );
  OR2_X1 U853 ( .A1(n799), .A2(n352), .ZN(n800) );
  NAND2_X1 U854 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U855 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U856 ( .A1(n804), .A2(n829), .ZN(n805) );
  XNOR2_X1 U857 ( .A(n806), .B(n805), .ZN(G75) );
  NAND2_X1 U858 ( .A1(G953), .A2(G224), .ZN(n807) );
  XNOR2_X1 U859 ( .A(KEYINPUT61), .B(n807), .ZN(n808) );
  NAND2_X1 U860 ( .A1(n808), .A2(G898), .ZN(n809) );
  NAND2_X1 U861 ( .A1(n810), .A2(n809), .ZN(n816) );
  XOR2_X1 U862 ( .A(G101), .B(n811), .Z(n813) );
  NOR2_X1 U863 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U864 ( .A(KEYINPUT125), .B(n814), .Z(n815) );
  XNOR2_X1 U865 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U866 ( .A(KEYINPUT124), .B(n817), .ZN(G69) );
  BUF_X1 U867 ( .A(n818), .Z(n819) );
  XNOR2_X1 U868 ( .A(n819), .B(n820), .ZN(n821) );
  XOR2_X1 U869 ( .A(n822), .B(n821), .Z(n828) );
  XOR2_X1 U870 ( .A(KEYINPUT126), .B(n828), .Z(n823) );
  XNOR2_X1 U871 ( .A(G227), .B(n823), .ZN(n824) );
  NAND2_X1 U872 ( .A1(n824), .A2(G900), .ZN(n825) );
  NAND2_X1 U873 ( .A1(n825), .A2(G953), .ZN(n832) );
  BUF_X1 U874 ( .A(n826), .Z(n827) );
  XNOR2_X1 U875 ( .A(n827), .B(n828), .ZN(n830) );
  NAND2_X1 U876 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U877 ( .A1(n832), .A2(n831), .ZN(G72) );
  XNOR2_X1 U878 ( .A(G137), .B(KEYINPUT127), .ZN(n834) );
  XNOR2_X1 U879 ( .A(n834), .B(n351), .ZN(G39) );
endmodule

