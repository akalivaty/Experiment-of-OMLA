//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT64), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n194), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  OAI211_X1 g018(.A(G128), .B(new_n201), .C1(new_n202), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n206), .B(new_n207), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .A3(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n212), .B1(new_n217), .B2(KEYINPUT3), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT73), .B(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(G101), .B1(new_n219), .B2(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT74), .B1(new_n219), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT74), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT75), .B1(new_n213), .B2(G104), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n211), .A3(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT10), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n199), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI211_X1 g048(.A(KEYINPUT76), .B(KEYINPUT10), .C1(new_n221), .C2(new_n231), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n212), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n214), .A2(G104), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G107), .ZN(new_n240));
  AOI21_X1  g054(.A(G107), .B1(new_n238), .B2(new_n239), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n237), .B(new_n240), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G101), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT0), .A4(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n202), .A2(new_n204), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(G101), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n220), .B(new_n237), .C1(new_n242), .C2(new_n241), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT4), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n233), .B2(new_n232), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n198), .B1(new_n236), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G101), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n228), .B1(new_n217), .B2(KEYINPUT74), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n224), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n237), .B1(new_n241), .B2(new_n242), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n240), .A2(new_n258), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n209), .B(new_n205), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n233), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT76), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n232), .A2(new_n199), .A3(new_n233), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n198), .ZN(new_n268));
  INV_X1    g082(.A(new_n232), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n269), .A2(KEYINPUT10), .B1(new_n251), .B2(new_n254), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n257), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n261), .A2(new_n262), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n210), .B1(new_n260), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g094(.A(KEYINPUT12), .B(new_n268), .C1(new_n280), .C2(new_n232), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n230), .A2(G101), .B1(new_n218), .B2(new_n220), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n205), .A2(new_n209), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n283), .A2(new_n284), .B1(new_n260), .B2(new_n263), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(new_n198), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n271), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n278), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G469), .B1(new_n289), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n287), .A2(new_n271), .A3(new_n277), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n236), .A2(new_n256), .A3(new_n198), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n268), .B1(new_n267), .B2(new_n270), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n276), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(new_n271), .A3(new_n277), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT77), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n292), .B(new_n293), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n277), .B1(new_n257), .B2(new_n271), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n300), .B1(new_n305), .B2(KEYINPUT77), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n294), .A2(new_n298), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT78), .A3(new_n292), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n291), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n211), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT69), .B1(new_n322), .B2(G146), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n319), .A2(new_n321), .A3(new_n324), .A4(new_n203), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n274), .A3(G214), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(KEYINPUT82), .B2(new_n200), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT82), .B(G143), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT18), .A3(G131), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT18), .A2(G131), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n331), .B(new_n335), .C1(new_n330), .C2(new_n332), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(G146), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n332), .A2(new_n330), .ZN(new_n343));
  NOR2_X1   g157(.A1(G237), .A2(G953), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n344), .A2(G214), .B1(new_n345), .B2(G143), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT17), .B(G131), .C1(new_n343), .C2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(KEYINPUT83), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n333), .A2(G131), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT17), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n331), .B(new_n351), .C1(new_n330), .C2(new_n332), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT83), .B1(new_n342), .B2(new_n347), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n317), .B(new_n337), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n349), .A2(new_n352), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n338), .A2(new_n339), .A3(G146), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n322), .B(KEYINPUT19), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(G146), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n337), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n317), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n315), .B1(new_n366), .B2(KEYINPUT20), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(KEYINPUT84), .A3(new_n368), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(KEYINPUT20), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n337), .B1(new_n354), .B2(new_n355), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n317), .ZN(new_n373));
  OAI21_X1  g187(.A(G475), .B1(new_n373), .B2(G902), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n274), .A2(G952), .ZN(new_n375));
  NAND2_X1  g189(.A1(G234), .A2(G237), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G902), .A3(G953), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT21), .B(G898), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G116), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G122), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n387), .A3(new_n213), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n208), .A2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n200), .A2(G128), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n389), .A2(new_n390), .B1(new_n393), .B2(new_n188), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n208), .A2(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n200), .A2(G128), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT13), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT85), .B1(new_n391), .B2(KEYINPUT13), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n394), .B1(new_n188), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n387), .A2(new_n406), .A3(KEYINPUT14), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n387), .B2(KEYINPUT14), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n385), .B1(new_n387), .B2(KEYINPUT14), .ZN(new_n411));
  OAI21_X1  g225(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n390), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n393), .A2(new_n188), .ZN(new_n414));
  OAI21_X1  g228(.A(G134), .B1(new_n391), .B2(new_n392), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n394), .B(KEYINPUT86), .C1(new_n188), .C2(new_n402), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n405), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G217), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n311), .A2(new_n420), .A3(G953), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n403), .A2(new_n404), .B1(new_n412), .B2(new_n416), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n418), .A3(new_n421), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n371), .A2(new_n374), .A3(new_n383), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n386), .A2(G119), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n434));
  INV_X1    g248(.A(G119), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(G116), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n386), .A2(KEYINPUT66), .A3(G119), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT5), .ZN(new_n439));
  INV_X1    g253(.A(G113), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT5), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(KEYINPUT2), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT2), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G113), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n439), .A2(new_n442), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n231), .A2(new_n447), .A3(new_n253), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n436), .A2(new_n437), .ZN(new_n451));
  INV_X1    g265(.A(new_n433), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n451), .A2(new_n452), .A3(new_n446), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n386), .A2(KEYINPUT66), .A3(G119), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT66), .B1(new_n386), .B2(G119), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n446), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n438), .A2(new_n446), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT67), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n245), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n448), .B1(new_n449), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n448), .B(new_n465), .C1(new_n449), .C2(new_n463), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n250), .A2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n284), .A2(new_n320), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G224), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n474), .B(KEYINPUT80), .Z(new_n475));
  XNOR2_X1  g289(.A(new_n472), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n465), .A2(KEYINPUT6), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n464), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n464), .B2(new_n478), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n469), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n283), .B(new_n447), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n465), .B(KEYINPUT8), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(new_n484), .B2(new_n474), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n474), .A2(new_n484), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n470), .A2(new_n471), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n482), .A2(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n488), .B2(new_n468), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n489), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n495), .A2(new_n494), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n432), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n314), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n435), .B2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(G119), .C2(new_n208), .ZN(new_n506));
  XNOR2_X1  g320(.A(G119), .B(G128), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  AOI22_X1  g322(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n341), .B2(new_n340), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n326), .A3(new_n358), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT22), .B(G137), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n512), .A3(new_n516), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n293), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n420), .B1(G234), .B2(new_n293), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT25), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(G902), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT71), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n530), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(KEYINPUT72), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n344), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n455), .A2(new_n462), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n193), .A2(new_n351), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n351), .B1(G134), .B2(new_n190), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n192), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n284), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n250), .A2(new_n198), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(KEYINPUT65), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n193), .A2(new_n351), .B1(new_n192), .B2(new_n543), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT65), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n284), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n541), .B1(new_n554), .B2(new_n547), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT28), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n249), .B1(new_n196), .B2(new_n197), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n551), .A2(new_n210), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT68), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n546), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n561), .A3(new_n541), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n540), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n547), .B2(new_n546), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n210), .B1(new_n545), .B2(KEYINPUT65), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n557), .B1(new_n568), .B2(new_n553), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(new_n566), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n548), .B(new_n540), .C1(new_n570), .C2(new_n541), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n547), .A2(new_n546), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT30), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n284), .B1(new_n552), .B2(new_n551), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n545), .A2(KEYINPUT65), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n566), .B(new_n547), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n541), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n549), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .A3(new_n540), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n565), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT32), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n556), .A2(new_n564), .ZN(new_n587));
  INV_X1    g401(.A(new_n540), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT31), .B1(new_n581), .B2(new_n540), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n541), .B1(new_n575), .B2(new_n578), .ZN(new_n591));
  NOR4_X1   g405(.A1(new_n591), .A2(new_n549), .A3(new_n572), .A4(new_n588), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n584), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n548), .B1(new_n570), .B2(new_n541), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n588), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT29), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n598), .B(new_n599), .C1(new_n587), .C2(new_n588), .ZN(new_n600));
  INV_X1    g414(.A(new_n564), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n580), .A2(new_n574), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n563), .B1(new_n602), .B2(new_n548), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n588), .A2(new_n599), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n536), .B1(new_n596), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n502), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  AND3_X1   g425(.A1(new_n481), .A2(new_n489), .A3(new_n491), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n491), .B1(new_n481), .B2(new_n489), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n497), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT89), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(KEYINPUT89), .B(new_n497), .C1(new_n612), .C2(new_n613), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n419), .A2(new_n422), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n421), .B1(new_n424), .B2(new_n418), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n423), .A2(new_n621), .A3(new_n425), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(G478), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n427), .A2(new_n293), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n426), .B2(new_n427), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n382), .B(new_n626), .C1(new_n371), .C2(new_n374), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n617), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT90), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT90), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n616), .A2(new_n630), .A3(new_n617), .A4(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n593), .B2(new_n293), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n583), .A2(new_n585), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n536), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n632), .A2(new_n314), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND2_X1   g454(.A1(new_n616), .A2(new_n617), .ZN(new_n641));
  INV_X1    g455(.A(new_n370), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n366), .A2(KEYINPUT20), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n374), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n382), .B(KEYINPUT91), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n644), .A2(new_n429), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n314), .A2(new_n641), .A3(new_n637), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n513), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n530), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n527), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n502), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(new_n655), .B1(new_n596), .B2(new_n608), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n616), .A3(new_n617), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n310), .A2(new_n661), .A3(new_n313), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n379), .A2(G900), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n377), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n644), .A2(new_n429), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(new_n664), .B(KEYINPUT39), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n314), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  INV_X1    g485(.A(new_n365), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n356), .B2(new_n363), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n369), .B1(new_n368), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT84), .B1(new_n673), .B2(new_n368), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n374), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n429), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n497), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n679), .A3(new_n654), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT94), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n602), .A2(new_n548), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n588), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT92), .ZN(new_n684));
  AOI21_X1  g498(.A(G902), .B1(new_n684), .B2(new_n571), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n596), .B1(new_n633), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT93), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n612), .A2(new_n613), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n498), .B1(new_n688), .B2(new_n494), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n681), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT95), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n671), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  INV_X1    g508(.A(new_n626), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n676), .A2(new_n695), .A3(new_n664), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n662), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  OAI21_X1  g513(.A(new_n293), .B1(new_n299), .B2(new_n301), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n313), .B1(new_n700), .B2(G469), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n306), .A2(new_n307), .ZN(new_n702));
  AND4_X1   g516(.A1(KEYINPUT78), .A2(new_n702), .A3(new_n292), .A4(new_n293), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT78), .B1(new_n308), .B2(new_n292), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n701), .B(new_n609), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n631), .B2(new_n629), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT41), .B(G113), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND3_X1  g522(.A1(new_n647), .A2(new_n616), .A3(new_n617), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND2_X1  g525(.A1(new_n432), .A2(new_n660), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n616), .A2(new_n617), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT96), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n312), .B1(new_n308), .B2(new_n292), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n304), .B2(new_n309), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT96), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n641), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n712), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n435), .ZN(G21));
  NAND4_X1  g535(.A1(new_n616), .A2(new_n676), .A3(new_n677), .A4(new_n617), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n584), .B(KEYINPUT97), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT98), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n601), .B2(new_n603), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n682), .A2(KEYINPUT28), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n728), .A3(new_n588), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n573), .A2(new_n582), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n634), .A2(new_n731), .A3(new_n532), .A4(new_n646), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n717), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND2_X1  g548(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n634), .A2(new_n731), .A3(new_n655), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT99), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n676), .A2(new_n737), .A3(new_n695), .A4(new_n664), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n715), .B2(new_n719), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT100), .B(G125), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G27));
  OAI21_X1  g556(.A(new_n290), .B1(new_n703), .B2(new_n704), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n735), .A2(new_n738), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n313), .A2(new_n679), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n689), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(new_n609), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n583), .A2(KEYINPUT32), .A3(new_n585), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n594), .B1(new_n593), .B2(new_n584), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n608), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n532), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT101), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n735), .A2(KEYINPUT42), .A3(new_n738), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n743), .A3(new_n747), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND4_X1  g577(.A1(new_n743), .A2(new_n609), .A3(new_n666), .A4(new_n747), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n304), .A2(new_n309), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n292), .B1(new_n289), .B2(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(KEYINPUT45), .B2(new_n289), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n772), .A2(KEYINPUT102), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(KEYINPUT102), .B2(new_n772), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n312), .ZN(new_n775));
  INV_X1    g589(.A(new_n676), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n695), .ZN(new_n777));
  NAND2_X1  g591(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n780));
  OAI21_X1  g594(.A(new_n779), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n636), .A3(new_n654), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n689), .A2(new_n679), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n775), .A2(new_n669), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT104), .B(G137), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G39));
  XOR2_X1   g605(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n792));
  NAND3_X1  g606(.A1(new_n774), .A2(new_n312), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n697), .A2(new_n536), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n787), .A2(new_n753), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT105), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n793), .B(new_n795), .C1(new_n775), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n781), .A2(new_n378), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n634), .A2(new_n731), .A3(new_n532), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n793), .B1(new_n775), .B2(new_n797), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n304), .A2(new_n309), .B1(G469), .B2(new_n700), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n313), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n787), .B(new_n804), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n690), .A2(new_n497), .A3(new_n713), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n803), .A3(new_n802), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT50), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n747), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT113), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n687), .A2(new_n536), .A3(new_n377), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n776), .A3(new_n626), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n736), .A3(new_n802), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(KEYINPUT50), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n812), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n800), .B(new_n801), .C1(new_n809), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n805), .A2(new_n808), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n804), .A2(new_n787), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n823), .B2(KEYINPUT112), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n759), .A3(new_n802), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n814), .A2(new_n676), .A3(new_n695), .A4(new_n815), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n713), .A2(KEYINPUT96), .A3(new_n714), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n718), .B1(new_n717), .B2(new_n641), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n803), .B(new_n802), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n375), .A3(new_n831), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT115), .B1(new_n827), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n820), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n701), .B(new_n732), .C1(new_n703), .C2(new_n704), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n709), .A2(new_n705), .B1(new_n839), .B2(new_n722), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n706), .ZN(new_n841));
  INV_X1    g655(.A(new_n712), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n829), .B2(new_n830), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n626), .B(new_n646), .C1(new_n371), .C2(new_n374), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n497), .A3(new_n499), .A4(new_n496), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT107), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT108), .B1(new_n676), .B2(new_n429), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT108), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n371), .A2(new_n677), .A3(new_n849), .A4(new_n374), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n689), .A3(new_n497), .A4(new_n645), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n689), .A2(KEYINPUT107), .A3(new_n497), .A4(new_n844), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n314), .A3(new_n637), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n314), .B(new_n501), .C1(new_n609), .C2(new_n656), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n841), .A2(new_n843), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n644), .A2(new_n677), .A3(new_n665), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n753), .A2(new_n654), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n739), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n743), .A3(new_n747), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n764), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n762), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n838), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n314), .A2(new_n641), .A3(new_n666), .A4(new_n660), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n740), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n655), .A2(new_n664), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT110), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n314), .A2(new_n686), .A3(new_n723), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n698), .A4(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n720), .A2(new_n706), .A3(new_n840), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n862), .B1(new_n750), .B2(new_n761), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n856), .A2(new_n855), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(KEYINPUT109), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n739), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n829), .B2(new_n830), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n667), .A3(new_n698), .A4(new_n871), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n865), .A2(new_n872), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n879), .B(new_n868), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT52), .B1(new_n866), .B2(new_n740), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n882), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n865), .A3(new_n876), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n837), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT111), .ZN(new_n889));
  INV_X1    g703(.A(new_n705), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n632), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n710), .A3(new_n733), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n892), .B2(new_n720), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT111), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n885), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n884), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n883), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n836), .A2(new_n888), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  INV_X1    g716(.A(new_n807), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(KEYINPUT49), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n754), .A2(new_n745), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n687), .A2(new_n690), .A3(new_n777), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT49), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n807), .B2(new_n907), .ZN(new_n908));
  OAI22_X1  g722(.A1(new_n901), .A2(new_n902), .B1(new_n904), .B2(new_n908), .ZN(G75));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n479), .A2(new_n480), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n469), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(new_n476), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  MUX2_X1   g729(.A(new_n910), .B(new_n911), .S(new_n915), .Z(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n293), .B1(new_n883), .B2(new_n898), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(G210), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n881), .A2(new_n882), .B1(new_n897), .B2(new_n884), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n920), .A2(KEYINPUT117), .A3(new_n921), .A4(new_n293), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n274), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n920), .A2(new_n921), .A3(new_n293), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n918), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT116), .B1(new_n930), .B2(new_n921), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n915), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n926), .A2(new_n932), .ZN(G51));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n920), .B2(new_n837), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n899), .A2(new_n934), .A3(KEYINPUT54), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n769), .B(KEYINPUT57), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n702), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n930), .A2(new_n768), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n924), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NAND2_X1  g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT120), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n930), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n925), .B1(new_n946), .B2(new_n364), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n364), .B2(new_n946), .ZN(G60));
  XOR2_X1   g762(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n624), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n900), .B2(new_n888), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n620), .A3(new_n622), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n620), .A2(new_n622), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n937), .A2(new_n953), .A3(new_n938), .A4(new_n950), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n954), .A3(new_n925), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n899), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n518), .A2(new_n519), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n899), .A2(new_n652), .A3(new_n957), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n925), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G66));
  NAND2_X1  g778(.A1(new_n857), .A2(new_n274), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT122), .Z(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n381), .B2(new_n473), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(G898), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n913), .B1(new_n969), .B2(G953), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n968), .B(new_n970), .Z(G69));
  XNOR2_X1  g785(.A(new_n570), .B(KEYINPUT123), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n359), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(G900), .B(G953), .C1(new_n974), .C2(G227), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(G227), .B2(new_n974), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n851), .B1(new_n676), .B2(new_n695), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n786), .A2(new_n609), .ZN(new_n978));
  OR3_X1    g792(.A1(new_n670), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n798), .A2(new_n789), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n867), .A2(new_n698), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n693), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n980), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n987), .B(new_n693), .C1(new_n982), .C2(new_n983), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n973), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n762), .A2(new_n798), .A3(new_n764), .A4(new_n789), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n774), .A2(new_n312), .A3(new_n669), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n759), .A2(new_n723), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT126), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n993), .A2(new_n984), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n998), .B2(new_n974), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n976), .B1(new_n992), .B2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(new_n597), .A2(new_n540), .ZN(new_n1001));
  INV_X1    g815(.A(new_n857), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n986), .B(new_n1002), .C1(new_n989), .C2(new_n990), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1001), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n883), .A2(new_n887), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n598), .A2(new_n571), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1007), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n993), .A2(new_n1002), .A3(new_n984), .A4(new_n997), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1010), .A2(new_n1005), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n581), .A2(new_n588), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n925), .B(new_n1009), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1006), .A2(new_n1014), .ZN(G57));
endmodule


