//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT39), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  OR2_X1    g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n207), .B2(new_n209), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(G155gat), .B2(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n208), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT69), .ZN(new_n225));
  INV_X1    g024(.A(G134gat), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n226), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G113gat), .A2(G120gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g029(.A1(G113gat), .A2(G120gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  AND2_X1   g034(.A1(G113gat), .A2(G120gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT70), .B1(new_n236), .B2(new_n228), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n230), .A4(new_n224), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n223), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n212), .B2(new_n239), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n233), .A2(new_n238), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT77), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n241), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n250), .A2(KEYINPUT84), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT84), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT77), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT77), .B1(new_n243), .B2(new_n245), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n240), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n251), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G1gat), .B(G29gat), .Z(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G57gat), .B(G85gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT84), .B1(new_n250), .B2(new_n251), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n256), .A2(new_n253), .A3(new_n257), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n221), .B(new_n239), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n202), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT40), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT5), .B1(new_n268), .B2(new_n251), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n240), .A2(new_n251), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n246), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n240), .A2(new_n279), .A3(new_n251), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n248), .B2(new_n249), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n264), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n259), .A2(KEYINPUT40), .A3(new_n265), .A4(new_n270), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n289), .A3(new_n293), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT65), .B1(new_n303), .B2(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n305), .B(new_n306), .C1(G169gat), .C2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT64), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT64), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n314), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT67), .B(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(G183gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n330), .B2(new_n319), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n326), .A2(new_n327), .B1(new_n314), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n328), .A2(new_n333), .A3(KEYINPUT28), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT28), .B1(new_n328), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n312), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n310), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n315), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n301), .B(new_n302), .C1(new_n332), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT67), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n329), .A2(KEYINPUT27), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G183gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n333), .A3(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT68), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n340), .A2(new_n342), .B1(G183gat), .B2(G190gat), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n302), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n331), .A2(new_n314), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n342), .A2(new_n304), .A3(new_n309), .A4(new_n307), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n324), .B1(new_n319), .B2(new_n321), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT64), .B(new_n320), .C1(new_n316), .C2(new_n318), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n369), .B2(KEYINPUT25), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n300), .B1(new_n346), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n326), .A2(new_n327), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n345), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT73), .B1(new_n374), .B2(new_n302), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n364), .C1(new_n332), .C2(new_n345), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n363), .B2(new_n370), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(new_n377), .C1(new_n364), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n299), .B(new_n380), .ZN(new_n381));
  AOI211_X1 g180(.A(new_n288), .B(new_n372), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT30), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n381), .ZN(new_n385));
  INV_X1    g184(.A(new_n372), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n287), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT74), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT68), .B1(new_n336), .B2(new_n344), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n301), .B1(new_n393), .B2(new_n332), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n364), .B1(new_n332), .B2(new_n345), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n302), .B1(new_n395), .B2(KEYINPUT73), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(new_n396), .B2(new_n377), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n288), .B1(new_n397), .B2(new_n372), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n385), .A2(KEYINPUT30), .A3(new_n386), .A4(new_n287), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n384), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n284), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n297), .B2(new_n298), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n222), .B1(new_n403), .B2(KEYINPUT80), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n212), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n223), .A2(new_n301), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n409), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n295), .B1(new_n293), .B2(new_n289), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n299), .B2(new_n413), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n221), .B1(new_n415), .B2(new_n222), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n299), .B1(new_n223), .B2(new_n301), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT81), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(KEYINPUT81), .A3(new_n418), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(G22gat), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  INV_X1    g222(.A(G50gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(KEYINPUT78), .B(KEYINPUT31), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G22gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n410), .A2(new_n418), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n428), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n410), .B2(new_n418), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT83), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n435), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n431), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n394), .A2(new_n302), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n443), .A2(new_n377), .A3(new_n375), .A4(new_n390), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n346), .A2(new_n371), .A3(new_n300), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n385), .A2(new_n386), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n288), .C1(new_n448), .C2(KEYINPUT37), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT38), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n448), .B2(KEYINPUT37), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n372), .B1(new_n379), .B2(new_n381), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n287), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n449), .A2(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n280), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n255), .B2(new_n254), .ZN(new_n457));
  OAI221_X1 g256(.A(KEYINPUT5), .B1(new_n251), .B2(new_n268), .C1(new_n275), .C2(new_n246), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n265), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n282), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT6), .B(new_n264), .C1(new_n278), .C2(new_n281), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n387), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n442), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n402), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n398), .A2(new_n399), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n383), .B1(new_n382), .B2(KEYINPUT30), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n387), .A2(KEYINPUT74), .A3(new_n388), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n442), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n244), .B1(new_n393), .B2(new_n332), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n370), .A2(new_n239), .A3(new_n391), .A4(new_n392), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  INV_X1    g274(.A(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n478), .B(KEYINPUT32), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n478), .B2(KEYINPUT32), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n479), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT71), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n474), .ZN(new_n489));
  INV_X1    g288(.A(new_n477), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT34), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n495), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n496), .A2(KEYINPUT36), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n472), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n496), .A2(new_n442), .A3(new_n498), .ZN(new_n503));
  INV_X1    g302(.A(new_n470), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n496), .A2(new_n442), .A3(new_n498), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n506), .A2(new_n470), .A3(KEYINPUT35), .ZN(new_n507));
  OAI22_X1  g306(.A1(new_n465), .A2(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g308(.A(new_n463), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n288), .B1(new_n448), .B2(KEYINPUT37), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT38), .B1(new_n452), .B2(new_n453), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT38), .B1(new_n454), .B2(new_n447), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n442), .C1(new_n284), .C2(new_n401), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n484), .A2(new_n485), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n497), .B1(new_n522), .B2(new_n483), .ZN(new_n523));
  INV_X1    g322(.A(new_n498), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n496), .A2(KEYINPUT36), .A3(new_n498), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(new_n527), .A3(new_n472), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT85), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n502), .A3(new_n504), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n506), .B2(new_n470), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n509), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT97), .ZN(new_n536));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  OR2_X1    g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G57gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G64gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(G64gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(KEYINPUT91), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n549), .A2(new_n545), .A3(G64gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G64gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT9), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n541), .A3(new_n542), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n558), .B(KEYINPUT7), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  OAI211_X1 g361(.A(G85gat), .B(G92gat), .C1(new_n562), .C2(KEYINPUT94), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G99gat), .B(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n564), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n557), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n540), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n556), .B1(new_n568), .B2(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n557), .A2(new_n570), .A3(KEYINPUT95), .A4(KEYINPUT10), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(new_n574), .ZN(new_n580));
  INV_X1    g379(.A(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n539), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n577), .B2(new_n578), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n577), .A2(new_n584), .A3(new_n578), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n538), .B1(new_n580), .B2(new_n581), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n586), .A2(KEYINPUT98), .A3(new_n587), .A4(new_n588), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n583), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(G29gat), .A2(G36gat), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n595), .A2(KEYINPUT14), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(KEYINPUT14), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT87), .B(G29gat), .ZN(new_n598));
  INV_X1    g397(.A(G36gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n602), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n604), .B(new_n605), .C1(new_n607), .C2(new_n600), .ZN(new_n608));
  INV_X1    g407(.A(new_n600), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n609), .A2(KEYINPUT88), .A3(new_n602), .A4(new_n606), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G15gat), .B(G22gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT16), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(G1gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(G1gat), .B2(new_n612), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G8gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n608), .A2(new_n610), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n615), .B(G8gat), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n608), .B2(new_n610), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n617), .B(new_n618), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT13), .Z(new_n634));
  NOR2_X1   g433(.A1(new_n611), .A2(new_n616), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n608), .A2(new_n610), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n624), .B2(new_n625), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n638), .B(new_n642), .C1(new_n624), .C2(new_n625), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT89), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n624), .A2(KEYINPUT89), .A3(new_n625), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n641), .A2(new_n643), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n632), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT92), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT93), .Z(new_n654));
  XOR2_X1   g453(.A(G134gat), .B(G162gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n623), .ZN(new_n658));
  INV_X1    g457(.A(new_n570), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n620), .A3(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n611), .A2(new_n570), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G190gat), .B(G218gat), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n657), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n656), .A3(new_n664), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G155gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G183gat), .B(G211gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT21), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n556), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(G127gat), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n621), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n682), .B2(new_n685), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n676), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n686), .A3(new_n675), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n594), .A2(new_n649), .A3(new_n671), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n534), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n468), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT99), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  INV_X1    g497(.A(new_n401), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n534), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT100), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT100), .B(new_n704), .C1(new_n700), .C2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n700), .A2(G8gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n705), .A4(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1325gat));
  OAI21_X1  g510(.A(G15gat), .B1(new_n695), .B2(new_n527), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n496), .A2(new_n498), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(G15gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n695), .B2(new_n714), .ZN(G1326gat));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n442), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  NOR3_X1   g517(.A1(new_n594), .A2(new_n649), .A3(new_n692), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n529), .B1(new_n528), .B2(new_n532), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n671), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n468), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(new_n598), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  INV_X1    g525(.A(new_n719), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n671), .B1(new_n720), .B2(new_n721), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n528), .A2(new_n532), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(KEYINPUT44), .A3(new_n670), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n727), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT102), .A3(new_n724), .ZN(new_n734));
  INV_X1    g533(.A(new_n598), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT102), .B1(new_n733), .B2(new_n724), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n722), .A2(G36gat), .A3(new_n401), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n731), .B1(KEYINPUT44), .B2(new_n728), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(new_n401), .A3(new_n727), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n599), .ZN(G1329gat));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n527), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n733), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n713), .A2(G43gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n751));
  INV_X1    g550(.A(new_n749), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n722), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n745), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n534), .B2(new_n671), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n747), .B(new_n719), .C1(new_n757), .C2(new_n731), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT47), .B1(new_n722), .B2(new_n752), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT105), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n763), .B(new_n760), .C1(new_n758), .C2(G43gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(G1330gat));
  NOR3_X1   g564(.A1(new_n722), .A2(G50gat), .A3(new_n442), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n742), .A2(new_n442), .A3(new_n727), .ZN(new_n769));
  OAI221_X1 g568(.A(new_n767), .B1(new_n768), .B2(KEYINPUT48), .C1(new_n769), .C2(new_n424), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n424), .B1(new_n733), .B2(new_n471), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n766), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1331gat));
  AOI22_X1  g573(.A1(new_n669), .A2(new_n667), .B1(new_n689), .B2(new_n691), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n594), .A2(new_n649), .A3(new_n775), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n730), .A2(KEYINPUT107), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT107), .B1(new_n730), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n468), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n545), .ZN(G1332gat));
  AOI21_X1  g580(.A(new_n401), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT108), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n779), .A2(KEYINPUT109), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT109), .B1(new_n779), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n552), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n784), .A2(new_n787), .A3(new_n552), .A4(new_n785), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n779), .B2(new_n527), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n713), .A2(G71gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n779), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1334gat));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n442), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(G78gat), .Z(G1335gat));
  INV_X1    g597(.A(new_n649), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n692), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n594), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n742), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n468), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n730), .A2(new_n670), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(KEYINPUT110), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n800), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n593), .A2(G85gat), .A3(new_n468), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT111), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n804), .A2(new_n815), .ZN(G1336gat));
  AOI21_X1  g615(.A(new_n560), .B1(new_n802), .B2(new_n699), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n401), .A2(G92gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n593), .B(new_n819), .C1(new_n808), .C2(new_n811), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n812), .A2(new_n594), .A3(new_n818), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n742), .A2(new_n401), .A3(new_n801), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n822), .B(new_n823), .C1(new_n560), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1337gat));
  OAI21_X1  g625(.A(G99gat), .B1(new_n803), .B2(new_n527), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n594), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n713), .A2(G99gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(G1338gat));
  INV_X1    g629(.A(G106gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n802), .B2(new_n471), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n442), .A2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n593), .B(new_n834), .C1(new_n808), .C2(new_n811), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT53), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n812), .A2(new_n594), .A3(new_n833), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n742), .A2(new_n442), .A3(new_n801), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n837), .B(new_n838), .C1(new_n831), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(G1339gat));
  NAND3_X1  g640(.A1(new_n649), .A2(new_n775), .A3(new_n593), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n591), .A2(new_n592), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(new_n587), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n573), .A2(new_n575), .A3(new_n581), .A4(new_n576), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT54), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n845), .A2(new_n585), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n538), .B1(new_n579), .B2(KEYINPUT54), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n849), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n586), .A2(new_n587), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT55), .B(new_n851), .C1(new_n852), .C2(new_n847), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n843), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n640), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n658), .A2(new_n621), .A3(new_n620), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n618), .B1(new_n856), .B2(new_n617), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n635), .A2(new_n637), .A3(new_n634), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n631), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n855), .A2(new_n669), .A3(new_n667), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n859), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n854), .A2(new_n649), .B1(new_n593), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n670), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n693), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT112), .B(new_n861), .C1(new_n863), .C2(new_n670), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n842), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n699), .A2(new_n468), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n503), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n799), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n870), .A2(KEYINPUT113), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(KEYINPUT113), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n799), .A2(G113gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n871), .B2(new_n594), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n594), .A2(G120gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(G1341gat));
  NAND4_X1  g679(.A1(new_n868), .A2(new_n503), .A3(new_n692), .A4(new_n869), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n681), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n693), .B1(new_n873), .B2(new_n874), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n681), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT115), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n884), .B(new_n888), .C1(new_n885), .C2(new_n681), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n671), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n670), .B1(new_n873), .B2(new_n874), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n226), .B2(new_n895), .ZN(G1343gat));
  NAND2_X1  g695(.A1(new_n869), .A2(new_n527), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n868), .B2(new_n471), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n670), .ZN(new_n901));
  INV_X1    g700(.A(new_n861), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n692), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n900), .B(new_n442), .C1(new_n904), .C2(new_n842), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n799), .B(new_n898), .C1(new_n899), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G141gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n649), .A2(G141gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n868), .A2(new_n471), .A3(new_n898), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT58), .B1(new_n906), .B2(G141gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n747), .A2(new_n468), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n868), .A2(new_n471), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT117), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n868), .A2(new_n917), .A3(new_n471), .A4(new_n914), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n916), .A2(new_n401), .A3(new_n908), .A4(new_n918), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n912), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n913), .B1(new_n912), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(G1344gat));
  NOR2_X1   g721(.A1(new_n593), .A2(G148gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n916), .A2(new_n401), .A3(new_n918), .A4(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n594), .B(new_n898), .C1(new_n899), .C2(new_n905), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT59), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT119), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n898), .A2(new_n594), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n842), .B(KEYINPUT121), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT122), .B1(new_n903), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n842), .B(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(new_n937), .C1(new_n692), .C2(new_n864), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n471), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n900), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n442), .A2(new_n900), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n868), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n932), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n926), .B1(new_n943), .B2(KEYINPUT123), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n939), .A2(new_n900), .B1(new_n868), .B2(new_n941), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n932), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n931), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n924), .B1(new_n930), .B2(new_n948), .ZN(G1345gat));
  OAI21_X1  g748(.A(new_n898), .B1(new_n899), .B2(new_n905), .ZN(new_n950));
  OAI21_X1  g749(.A(G155gat), .B1(new_n950), .B2(new_n693), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n693), .A2(G155gat), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n916), .A2(new_n401), .A3(new_n918), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1346gat));
  INV_X1    g753(.A(new_n950), .ZN(new_n955));
  INV_X1    g754(.A(G162gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n670), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n916), .A2(new_n401), .A3(new_n671), .A4(new_n918), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n955), .A2(new_n957), .B1(new_n958), .B2(new_n956), .ZN(G1347gat));
  AND2_X1   g758(.A1(new_n868), .A2(new_n503), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n401), .A2(new_n724), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(G169gat), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(new_n649), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n962), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n799), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n964), .B1(new_n967), .B2(new_n963), .ZN(G1348gat));
  INV_X1    g767(.A(G176gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n969), .A3(new_n594), .ZN(new_n970));
  OAI21_X1  g769(.A(G176gat), .B1(new_n962), .B2(new_n593), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1349gat));
  OR3_X1    g771(.A1(new_n962), .A2(new_n333), .A3(new_n693), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n329), .B1(new_n962), .B2(new_n693), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n973), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n966), .A2(new_n328), .A3(new_n671), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n671), .A3(new_n961), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n982));
  AND4_X1   g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(G190gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n347), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n981), .A2(new_n984), .B1(new_n980), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n979), .B1(new_n983), .B2(new_n985), .ZN(G1351gat));
  INV_X1    g785(.A(new_n961), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n747), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n946), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n649), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AND4_X1   g791(.A1(new_n471), .A2(new_n868), .A3(new_n527), .A4(new_n961), .ZN(new_n993));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n799), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n946), .A2(new_n989), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n994), .B1(new_n997), .B2(new_n799), .ZN(new_n998));
  INV_X1    g797(.A(new_n995), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT126), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n996), .A2(new_n1000), .ZN(G1352gat));
  INV_X1    g800(.A(G204gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n993), .A2(new_n1002), .A3(new_n594), .ZN(new_n1003));
  XOR2_X1   g802(.A(new_n1003), .B(KEYINPUT62), .Z(new_n1004));
  OAI21_X1  g803(.A(G204gat), .B1(new_n990), .B2(new_n593), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1353gat));
  NAND3_X1  g805(.A1(new_n993), .A2(new_n291), .A3(new_n692), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n997), .A2(new_n692), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(G1354gat));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n671), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(new_n292), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n997), .A2(G218gat), .A3(new_n671), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(G1355gat));
endmodule


