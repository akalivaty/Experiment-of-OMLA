//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT76), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(G211gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(G211gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT75), .B(G211gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT22), .B1(new_n212), .B2(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(G204gat), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(G197gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(G204gat), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n211), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n226));
  OAI21_X1  g025(.A(G218gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n229), .A2(new_n210), .A3(new_n222), .A4(new_n217), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT3), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT2), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n237), .B2(KEYINPUT2), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G141gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G141gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n245), .A2(new_n247), .A3(G148gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n244), .B2(G148gat), .ZN(new_n250));
  INV_X1    g049(.A(G148gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT81), .B1(new_n251), .B2(G141gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(new_n247), .A3(G148gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n243), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n244), .A2(G148gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n251), .A2(G141gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n236), .A2(KEYINPUT79), .A3(new_n237), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n205), .B1(new_n233), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n243), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT82), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n269), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n231), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n231), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n261), .A2(KEYINPUT3), .A3(new_n270), .ZN(new_n283));
  INV_X1    g082(.A(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n269), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n224), .B2(new_n230), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(KEYINPUT3), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n285), .A2(KEYINPUT87), .A3(new_n205), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G22gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n229), .A2(new_n222), .A3(new_n217), .ZN(new_n292));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n284), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n293), .B2(new_n292), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n271), .B1(new_n295), .B2(new_n277), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n280), .A2(new_n296), .B1(new_n203), .B2(new_n204), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G78gat), .B(G106gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT86), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G50gat), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n291), .B1(new_n290), .B2(new_n297), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n304), .A2(KEYINPUT90), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT90), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT88), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n290), .A2(KEYINPUT88), .A3(new_n291), .A4(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n297), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G22gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315));
  INV_X1    g114(.A(new_n303), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n308), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OR3_X1    g124(.A1(new_n323), .A2(KEYINPUT26), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT28), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n323), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n327), .A2(new_n328), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n326), .A2(new_n331), .A3(new_n332), .A4(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n322), .B2(KEYINPUT23), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT24), .ZN(new_n346));
  INV_X1    g145(.A(G183gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(new_n328), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT64), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n328), .A3(KEYINPUT65), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT64), .B(new_n346), .C1(new_n347), .C2(new_n328), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT25), .B1(new_n345), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n348), .B(new_n356), .C1(G183gat), .C2(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n343), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n325), .B1(KEYINPUT23), .B2(new_n322), .ZN(new_n361));
  AND4_X1   g160(.A1(KEYINPUT25), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n336), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n363), .A2(new_n232), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n231), .B(new_n365), .C1(new_n366), .C2(new_n364), .ZN(new_n367));
  INV_X1    g166(.A(new_n365), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n363), .B2(new_n279), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n282), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n370), .A3(new_n374), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT30), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G127gat), .B(G134gat), .Z(new_n381));
  OR2_X1    g180(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n381), .B(new_n382), .C1(KEYINPUT1), .C2(new_n384), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT84), .B1(new_n271), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391));
  NOR4_X1   g190(.A1(new_n261), .A2(new_n390), .A3(new_n270), .A4(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT4), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n276), .A2(new_n388), .A3(new_n269), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n261), .B2(new_n270), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n278), .A2(new_n398), .A3(new_n390), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n391), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n271), .A2(KEYINPUT84), .A3(new_n388), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n286), .A2(new_n390), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n401), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n404), .A3(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n401), .A3(new_n399), .A4(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n397), .A2(new_n402), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  AOI21_X1  g215(.A(KEYINPUT6), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n416), .B2(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n411), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n393), .A3(new_n396), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n416), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n380), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n308), .B(KEYINPUT91), .C1(new_n317), .C2(new_n318), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n321), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n416), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n412), .A2(KEYINPUT92), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n432), .B2(new_n417), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n375), .B1(new_n371), .B2(KEYINPUT37), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n282), .B(new_n365), .C1(new_n366), .C2(new_n364), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n231), .B1(new_n368), .B2(new_n369), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT37), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n378), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n367), .B2(new_n370), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT38), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT93), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT93), .B(KEYINPUT38), .C1(new_n434), .C2(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n393), .A2(new_n399), .A3(new_n396), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n407), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n448), .A2(new_n407), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT39), .B1(new_n406), .B2(new_n407), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n416), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n454), .A2(KEYINPUT40), .B1(new_n430), .B2(new_n431), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n377), .A2(new_n379), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n433), .A2(new_n447), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n363), .A2(new_n390), .ZN(new_n459));
  AND2_X1   g258(.A1(G227gat), .A2(G233gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n388), .B(new_n336), .C1(new_n358), .C2(new_n362), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT34), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n459), .A2(new_n462), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT32), .B1(new_n466), .B2(new_n461), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n461), .B1(new_n459), .B2(new_n462), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n470), .ZN(new_n477));
  INV_X1    g276(.A(new_n471), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT71), .B1(new_n474), .B2(new_n475), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n473), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n465), .B1(new_n482), .B2(KEYINPUT72), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n467), .A2(new_n472), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(KEYINPUT32), .C1(new_n466), .C2(new_n461), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n471), .B1(new_n466), .B2(new_n461), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n481), .A4(new_n477), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT72), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n464), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n484), .A2(new_n488), .A3(new_n464), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n464), .B1(new_n484), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n492), .A2(KEYINPUT36), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n458), .A2(new_n319), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n319), .A2(new_n424), .A3(new_n492), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n494), .A2(new_n495), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n504), .A2(KEYINPUT35), .A3(new_n380), .ZN(new_n505));
  INV_X1    g304(.A(new_n433), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n319), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n427), .A2(new_n500), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT14), .B(G29gat), .Z(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G36gat), .ZN(new_n512));
  INV_X1    g311(.A(G43gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(G50gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n512), .B1(KEYINPUT15), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(G50gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(KEYINPUT15), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(KEYINPUT15), .A3(new_n519), .A4(new_n518), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT95), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n528), .A2(KEYINPUT95), .A3(G1gat), .ZN(new_n531));
  OAI221_X1 g330(.A(new_n526), .B1(G1gat), .B2(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n521), .A2(new_n522), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n534), .B(new_n535), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n538), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n542), .A2(new_n552), .A3(new_n546), .A4(new_n543), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g358(.A(G71gat), .ZN(new_n560));
  INV_X1    g359(.A(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G127gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n534), .B1(new_n566), .B2(new_n565), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n234), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n570), .A2(new_n571), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n571), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT97), .Z(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n587), .B2(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n596), .A3(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n525), .A2(new_n536), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT99), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n600), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n523), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n603), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n586), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n585), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n608), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n204), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n565), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  INV_X1    g421(.A(new_n564), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n563), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n598), .A3(new_n599), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n625), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(new_n620), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  OR2_X1    g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n582), .A2(new_n618), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n508), .A2(new_n557), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n418), .A2(new_n423), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n380), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT42), .ZN(new_n646));
  INV_X1    g445(.A(new_n639), .ZN(new_n647));
  INV_X1    g446(.A(new_n380), .ZN(new_n648));
  OAI21_X1  g447(.A(G8gat), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT101), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(G8gat), .C1(new_n647), .C2(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n646), .A2(new_n655), .A3(new_n650), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n498), .A2(new_n499), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n647), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n504), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n647), .B2(new_n660), .ZN(G1326gat));
  AND2_X1   g460(.A1(new_n321), .A2(new_n426), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NOR2_X1   g464(.A1(new_n508), .A2(new_n557), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n582), .A2(new_n618), .A3(new_n636), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n509), .A3(new_n641), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT44), .B1(new_n508), .B2(new_n618), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n500), .A2(new_n427), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n502), .A2(new_n507), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT104), .B1(new_n614), .B2(new_n617), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n613), .A2(new_n611), .A3(new_n609), .ZN(new_n677));
  INV_X1    g476(.A(new_n586), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n616), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n672), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n582), .B(KEYINPUT103), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n557), .A3(new_n636), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n640), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(new_n689), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n380), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n689), .B2(new_n648), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(G36gat), .A3(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n668), .A2(G36gat), .A3(new_n648), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1329gat));
  OAI21_X1  g498(.A(G43gat), .B1(new_n689), .B2(new_n658), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n669), .A2(new_n513), .A3(new_n503), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT47), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n702), .B(new_n704), .ZN(G1330gat));
  INV_X1    g504(.A(new_n515), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n669), .A2(new_n662), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n662), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n515), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n319), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n706), .B1(new_n692), .B2(new_n712), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n709), .A2(KEYINPUT48), .B1(new_n711), .B2(new_n713), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n582), .A2(new_n618), .A3(new_n557), .A4(new_n636), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n508), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n641), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n380), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  INV_X1    g521(.A(new_n658), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n560), .B1(new_n716), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n504), .A2(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n662), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n582), .A2(new_n556), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n637), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n672), .B2(new_n684), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n640), .ZN(new_n736));
  INV_X1    g535(.A(new_n618), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n675), .A2(new_n737), .A3(new_n730), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n737), .A4(new_n730), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT107), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n641), .A2(new_n587), .A3(new_n636), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n736), .B1(new_n743), .B2(new_n744), .ZN(G1336gat));
  AOI21_X1  g544(.A(new_n588), .B1(new_n734), .B2(new_n380), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n648), .A2(new_n637), .A3(G92gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n740), .B2(new_n741), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n675), .B2(new_n737), .ZN(new_n753));
  INV_X1    g552(.A(new_n683), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n508), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n380), .B(new_n732), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G92gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n751), .B1(new_n757), .B2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n747), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n750), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n750), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1337gat));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n735), .B2(new_n658), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n734), .A2(KEYINPUT110), .A3(new_n723), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(G99gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n504), .A2(G99gat), .A3(new_n637), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT111), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n743), .B2(new_n770), .ZN(G1338gat));
  INV_X1    g570(.A(G106gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n734), .B2(new_n662), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n712), .A2(new_n772), .A3(new_n636), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n773), .B1(new_n742), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n772), .B1(new_n734), .B2(new_n712), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n742), .A2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n777), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n780), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n638), .A2(new_n556), .ZN(new_n782));
  INV_X1    g581(.A(new_n628), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n626), .A2(new_n627), .A3(new_n620), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n633), .B1(new_n628), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n789), .B(new_n633), .C1(new_n628), .C2(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(KEYINPUT55), .B(new_n785), .C1(new_n788), .C2(new_n790), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n556), .A3(new_n635), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n544), .A2(new_n545), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n551), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n555), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n636), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n682), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n614), .A2(KEYINPUT104), .A3(new_n617), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n680), .B1(new_n679), .B2(new_n616), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n793), .A2(new_n799), .A3(new_n635), .A4(new_n794), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n782), .B1(new_n809), .B2(new_n686), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n640), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n319), .A2(new_n492), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n648), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT113), .Z(new_n815));
  INV_X1    g614(.A(G113gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n556), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n810), .A2(new_n662), .A3(new_n504), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n640), .A2(new_n380), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n557), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n823), .A3(new_n636), .ZN(new_n824));
  OAI21_X1  g623(.A(G120gat), .B1(new_n820), .B2(new_n637), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1341gat));
  INV_X1    g625(.A(new_n582), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n814), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(G127gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n818), .A2(G127gat), .A3(new_n687), .A4(new_n819), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n618), .A2(new_n380), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n813), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n820), .B2(new_n618), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n682), .A2(new_n806), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n795), .A2(new_n800), .B1(new_n676), .B2(new_n681), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n686), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n782), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n319), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(KEYINPUT57), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT115), .B(new_n847), .C1(new_n810), .C2(new_n319), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n849));
  NAND2_X1  g648(.A1(new_n791), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n556), .A3(new_n635), .A4(new_n794), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n800), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n851), .B2(new_n800), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n618), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n808), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n782), .B1(new_n857), .B2(new_n827), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n662), .A2(KEYINPUT57), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n846), .B(new_n848), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n658), .A2(new_n819), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n556), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n245), .A2(new_n247), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n723), .A2(new_n319), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n811), .A2(new_n866), .ZN(new_n867));
  AND4_X1   g666(.A1(new_n244), .A2(new_n867), .A3(new_n648), .A4(new_n556), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n863), .A2(new_n871), .A3(new_n864), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n863), .B2(new_n864), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  AND2_X1   g675(.A1(new_n867), .A2(new_n648), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n251), .A3(new_n636), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n862), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n637), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(KEYINPUT59), .A3(new_n251), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n851), .A2(new_n800), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n737), .B1(new_n883), .B2(new_n853), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n806), .A2(new_n618), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n827), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n844), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n847), .A3(new_n662), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n810), .B2(new_n319), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n636), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G148gat), .B1(new_n890), .B2(new_n861), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n878), .B1(new_n881), .B2(new_n892), .ZN(G1345gat));
  OAI21_X1  g692(.A(G155gat), .B1(new_n879), .B2(new_n686), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n234), .A3(new_n582), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n879), .B2(new_n682), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n235), .A3(new_n835), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n641), .A2(new_n648), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n818), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n557), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT121), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n810), .A2(new_n641), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(new_n380), .A3(new_n812), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n337), .A3(new_n556), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n338), .A3(new_n636), .ZN(new_n910));
  OAI21_X1  g709(.A(G176gat), .B1(new_n903), .B2(new_n637), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT122), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n327), .A3(new_n582), .ZN(new_n914));
  OAI21_X1  g713(.A(G183gat), .B1(new_n903), .B2(new_n686), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n907), .A2(new_n328), .A3(new_n805), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT124), .ZN(new_n920));
  OAI21_X1  g719(.A(G190gat), .B1(new_n903), .B2(new_n618), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(G1351gat));
  AND3_X1   g724(.A1(new_n906), .A2(new_n380), .A3(new_n866), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n556), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n658), .A2(new_n902), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n888), .A2(new_n889), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n557), .A2(new_n219), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n637), .A2(G204gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n890), .B2(new_n928), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1353gat));
  INV_X1    g742(.A(new_n212), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n944), .A3(new_n582), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n888), .A2(new_n582), .A3(new_n889), .A4(new_n929), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n926), .A2(new_n207), .A3(new_n805), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(new_n618), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n207), .ZN(G1355gat));
endmodule


