//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  INV_X1    g0008(.A(G264), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n201), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT66), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT0), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n227), .A2(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n233), .B1(new_n232), .B2(new_n231), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n220), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G97), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n226), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n222), .B2(new_n224), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT8), .B(G58), .Z(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n255), .A2(new_n256), .B1(G150), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT71), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n253), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT72), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n268), .A2(new_n265), .A3(G13), .A4(G20), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n264), .B1(new_n270), .B2(new_n253), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(G20), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n253), .B1(new_n267), .B2(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n271), .A2(G50), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n263), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT69), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n287), .A2(new_n292), .A3(G222), .A4(new_n288), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT68), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT68), .B1(new_n284), .B2(new_n285), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G77), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT70), .B(G223), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n287), .A2(G1698), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n291), .A2(new_n293), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(G274), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n310), .B2(G226), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n278), .B1(new_n312), .B2(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(new_n311), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n278), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n312), .A2(G190), .B1(KEYINPUT9), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n314), .A2(G200), .B1(new_n278), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n323), .A3(new_n320), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n316), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n308), .B1(new_n310), .B2(G238), .ZN(new_n327));
  INV_X1    g0127(.A(G97), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n254), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G226), .A2(G1698), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n207), .B2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n287), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n327), .B1(new_n332), .B2(new_n302), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n327), .B(new_n335), .C1(new_n332), .C2(new_n302), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n326), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(G179), .A3(new_n336), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n255), .ZN(new_n343));
  INV_X1    g0143(.A(G77), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n257), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n346), .A2(new_n276), .B1(new_n221), .B2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n253), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT11), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n270), .A2(new_n202), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n273), .A2(G68), .A3(new_n272), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n334), .A2(new_n336), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(G200), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n334), .A2(KEYINPUT74), .A3(G190), .A4(new_n336), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n256), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n225), .A2(new_n344), .B1(new_n363), .B2(new_n346), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n343), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n253), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n273), .A2(G77), .A3(new_n272), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n267), .A2(new_n269), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(G77), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n371), .B1(new_n208), .B2(new_n287), .C1(new_n289), .C2(new_n207), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n303), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n308), .B1(new_n310), .B2(G244), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n376), .B2(G190), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n370), .B1(new_n376), .B2(G169), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G179), .B2(new_n375), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n325), .A2(new_n362), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT18), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n272), .B1(new_n273), .B2(KEYINPUT73), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n264), .B(new_n253), .C1(new_n267), .C2(new_n269), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n386), .A2(new_n387), .A3(new_n363), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n369), .A2(new_n256), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n271), .A2(new_n272), .A3(new_n256), .A4(new_n274), .ZN(new_n391));
  INV_X1    g0191(.A(new_n389), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(KEYINPUT75), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n283), .A2(new_n395), .A3(new_n221), .A4(new_n286), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n222), .A2(new_n224), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT3), .B(G33), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT7), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n396), .A2(G68), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(G159), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(new_n346), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n394), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n401), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n284), .B2(new_n285), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n407), .B2(new_n395), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n284), .A2(new_n285), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n225), .A2(new_n409), .A3(new_n395), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT16), .B(new_n406), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n411), .A2(new_n253), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n390), .A2(new_n393), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n284), .A2(new_n285), .A3(G223), .A4(new_n288), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  INV_X1    g0215(.A(G87), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n254), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(G226), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n398), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n398), .A2(new_n420), .A3(G223), .A4(new_n288), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n415), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n303), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n307), .B1(new_n207), .B2(new_n309), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT77), .B1(new_n426), .B2(G179), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n422), .B2(new_n303), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n326), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n384), .B1(new_n413), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n405), .A2(new_n412), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n388), .A2(new_n385), .A3(new_n389), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT75), .B1(new_n391), .B2(new_n392), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n428), .A2(G169), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n378), .B1(new_n423), .B2(new_n425), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n359), .B(new_n424), .C1(new_n422), .C2(new_n303), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n435), .C1(new_n436), .C2(new_n437), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT17), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n413), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n383), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT79), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n369), .A2(new_n328), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n265), .A2(G33), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n273), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n458), .B(new_n459), .C1(new_n462), .C2(new_n328), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n328), .B1(new_n273), .B2(new_n460), .ZN(new_n464));
  INV_X1    g0264(.A(new_n459), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT79), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n208), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  INV_X1    g0268(.A(new_n249), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(KEYINPUT6), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(new_n397), .B1(G77), .B2(new_n257), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n396), .A2(G107), .A3(new_n399), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n253), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  INV_X1    g0276(.A(G244), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n288), .B(new_n478), .C1(new_n294), .C2(new_n295), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n284), .A2(new_n285), .A3(G244), .A4(new_n288), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(new_n476), .B1(G33), .B2(G283), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n303), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G41), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n265), .A2(G45), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(new_n302), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  INV_X1    g0292(.A(new_n490), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(G274), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(KEYINPUT80), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n378), .B1(new_n484), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n359), .B(new_n495), .C1(new_n483), .C2(new_n303), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n475), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n484), .A2(new_n430), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n495), .B1(new_n483), .B2(new_n303), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(G169), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n463), .A2(new_n466), .B1(new_n473), .B2(new_n253), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT81), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n326), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT81), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n475), .A3(new_n510), .A4(new_n503), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n502), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n303), .B1(new_n493), .B2(new_n492), .ZN(new_n513));
  INV_X1    g0313(.A(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G250), .B2(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n409), .B1(new_n254), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(G264), .A2(new_n513), .B1(new_n518), .B2(new_n303), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(KEYINPUT85), .A3(new_n359), .A4(new_n494), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  OAI211_X1 g0321(.A(G264), .B(new_n302), .C1(new_n489), .C2(new_n490), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n514), .B2(G1698), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n398), .B1(G33), .B2(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n494), .B(new_n522), .C1(new_n525), .C2(new_n302), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n521), .B1(new_n526), .B2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n378), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT23), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT82), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n531), .B(new_n533), .C1(new_n221), .C2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n222), .A2(new_n224), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n225), .A2(new_n398), .A3(KEYINPUT22), .A4(G87), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n416), .B1(new_n283), .B2(new_n286), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n296), .B2(new_n416), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT24), .A3(new_n539), .A4(new_n538), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(new_n253), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n369), .B2(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n208), .B2(new_n461), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n529), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n526), .A2(new_n556), .A3(G169), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n556), .B1(new_n526), .B2(G169), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n526), .A2(new_n430), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n253), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n541), .B2(new_n542), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n552), .B1(new_n563), .B2(new_n546), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n555), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n547), .A2(new_n553), .ZN(new_n566));
  INV_X1    g0366(.A(new_n559), .ZN(new_n567));
  INV_X1    g0367(.A(new_n560), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n557), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(KEYINPUT84), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n554), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n416), .A2(new_n328), .A3(new_n208), .ZN(new_n572));
  AND3_X1   g0372(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n397), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n225), .A2(new_n398), .A3(G68), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT19), .B1(new_n255), .B2(G97), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n253), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n462), .A2(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n270), .A2(new_n365), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n302), .A2(G250), .A3(new_n490), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n493), .A2(G274), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G238), .A2(G1698), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n477), .B2(G1698), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(new_n398), .B1(G33), .B2(G116), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n302), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n584), .B(G190), .C1(new_n302), .C2(new_n587), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n398), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G116), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n302), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n582), .A2(new_n583), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n326), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n584), .B(new_n430), .C1(new_n302), .C2(new_n587), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n365), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n462), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n578), .A2(new_n600), .A3(new_n580), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n581), .A2(new_n591), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G283), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n225), .B(new_n603), .C1(G33), .C2(new_n328), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n252), .A2(new_n226), .B1(G20), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT20), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n328), .B2(G33), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT20), .B(new_n606), .C1(new_n397), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n273), .A2(G116), .A3(new_n460), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G116), .B2(new_n369), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n283), .A2(G303), .A3(new_n286), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n209), .A2(G1698), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n398), .B(new_n616), .C1(G257), .C2(G1698), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n302), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n302), .B1(new_n489), .B2(new_n490), .ZN(new_n619));
  INV_X1    g0419(.A(G270), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n494), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n614), .B1(new_n378), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(G190), .B2(new_n622), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  OAI21_X1  g0425(.A(G169), .B1(new_n618), .B2(new_n621), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n614), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n626), .ZN(new_n628));
  OAI221_X1 g0428(.A(new_n612), .B1(G116), .B2(new_n369), .C1(new_n607), .C2(new_n610), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(KEYINPUT21), .A3(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n618), .A2(new_n430), .A3(new_n621), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n512), .A2(new_n571), .A3(new_n602), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n457), .A2(new_n635), .ZN(G372));
  AOI21_X1  g0436(.A(new_n380), .B1(new_n430), .B2(new_n376), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n361), .B1(new_n342), .B2(new_n353), .ZN(new_n638));
  INV_X1    g0438(.A(new_n452), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n444), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n322), .A2(new_n324), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n316), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n303), .A2(new_n483), .B1(new_n497), .B2(new_n498), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n508), .A2(new_n326), .B1(new_n643), .B2(new_n430), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n602), .A2(new_n644), .A3(new_n645), .A4(new_n475), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n598), .A2(new_n601), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n507), .A2(new_n602), .A3(new_n511), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(KEYINPUT26), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n633), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n566), .A2(new_n569), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n554), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n512), .A2(new_n653), .A3(new_n602), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n642), .B1(new_n457), .B2(new_n657), .ZN(G369));
  OR2_X1    g0458(.A1(new_n634), .A2(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n634), .A2(KEYINPUT86), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n225), .A2(G13), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n265), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n659), .B(new_n660), .C1(new_n614), .C2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n614), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n633), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n652), .A2(new_n668), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n566), .A2(new_n667), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n571), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n571), .A2(new_n633), .A3(new_n668), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n667), .B(KEYINPUT87), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n652), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n230), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n572), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n228), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n522), .B1(new_n525), .B2(new_n302), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n588), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n504), .A2(new_n631), .A3(KEYINPUT30), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT88), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n504), .A2(new_n631), .A3(new_n694), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n526), .A2(new_n588), .A3(new_n430), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n643), .A2(new_n622), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT88), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n667), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n699), .A3(new_n695), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n682), .A2(new_n708), .A3(KEYINPUT31), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n709), .C1(new_n635), .C2(new_n682), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(KEYINPUT89), .A3(G330), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n561), .A2(new_n564), .A3(new_n555), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT84), .B1(new_n566), .B2(new_n569), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n651), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n512), .A3(new_n602), .A4(new_n654), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n505), .A2(new_n506), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT26), .A3(new_n602), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT90), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT90), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n720), .A2(new_n723), .A3(KEYINPUT26), .A4(new_n602), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n649), .A2(new_n645), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n719), .B(new_n647), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n668), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n682), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n656), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  OR4_X1    g0532(.A1(KEYINPUT91), .A2(new_n715), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n729), .A2(new_n732), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT91), .B1(new_n734), .B2(new_n715), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n692), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n265), .B1(new_n661), .B2(G45), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n688), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT92), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n287), .A2(G355), .A3(new_n230), .ZN(new_n743));
  INV_X1    g0543(.A(G45), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n247), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n686), .A2(new_n398), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G45), .B2(new_n228), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n743), .B1(G116), .B2(new_n230), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n226), .B1(G20), .B2(new_n326), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n742), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n359), .A2(new_n378), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n397), .A2(G179), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G326), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n359), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n225), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n225), .A2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n430), .A2(G200), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n760), .B1(new_n517), .B2(new_n762), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT94), .Z(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n430), .A3(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n763), .A2(new_n430), .A3(new_n378), .ZN(new_n772));
  INV_X1    g0572(.A(G329), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n757), .A2(G20), .A3(new_n430), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n225), .A2(new_n430), .A3(new_n359), .A4(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n296), .B1(new_n775), .B2(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n763), .A2(G179), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n774), .B(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n776), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n296), .B1(G87), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n762), .A2(new_n328), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n208), .C2(new_n771), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n766), .A2(new_n344), .B1(new_n202), .B2(new_n781), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n778), .A2(new_n201), .B1(new_n276), .B2(new_n758), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n772), .A2(new_n403), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n769), .A2(new_n784), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n752), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n755), .B1(new_n756), .B2(new_n795), .C1(new_n672), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n742), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n675), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n672), .A2(G330), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(G396));
  AOI22_X1  g0602(.A1(new_n765), .A2(G159), .B1(G143), .B2(new_n777), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  INV_X1    g0604(.A(G150), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(new_n804), .B2(new_n758), .C1(new_n805), .C2(new_n781), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT34), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n398), .B1(new_n776), .B2(new_n276), .C1(new_n762), .C2(new_n201), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n771), .A2(new_n202), .ZN(new_n811));
  INV_X1    g0611(.A(new_n772), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n811), .C1(G132), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n296), .B1(new_n208), .B2(new_n776), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n787), .B(new_n815), .C1(G311), .C2(new_n812), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n759), .A2(G303), .B1(new_n777), .B2(G294), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n782), .A2(G283), .B1(new_n765), .B2(G116), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n771), .A2(new_n416), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n821), .A2(KEYINPUT95), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n753), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n753), .A2(new_n749), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n798), .C1(G77), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  NAND2_X1  g0629(.A1(new_n667), .A2(new_n370), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n637), .B1(new_n379), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n382), .A2(new_n667), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n751), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT97), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n715), .B(new_n833), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(new_n731), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n798), .B1(new_n836), .B2(new_n731), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  OR2_X1    g0640(.A1(new_n705), .A2(new_n706), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n707), .C1(new_n635), .C2(new_n682), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n456), .A2(G330), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n353), .B(new_n667), .C1(new_n339), .C2(new_n341), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT98), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n353), .A2(new_n667), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n354), .A2(new_n361), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n842), .A2(new_n849), .A3(new_n833), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n434), .A2(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n411), .A2(new_n253), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n225), .A2(new_n409), .A3(new_n395), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n853), .B(G68), .C1(new_n395), .C2(new_n407), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n854), .B2(new_n406), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n392), .B(new_n391), .C1(new_n852), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n665), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT100), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n431), .A3(new_n427), .A4(new_n432), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n448), .A2(new_n860), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT101), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT37), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n438), .B1(new_n442), .B2(new_n857), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(new_n448), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT100), .ZN(new_n870));
  INV_X1    g0670(.A(new_n858), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n453), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n859), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n859), .A2(new_n869), .A3(new_n872), .A4(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n850), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n413), .B1(new_n433), .B2(new_n665), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n880), .B2(KEYINPUT102), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT103), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n866), .A2(new_n882), .A3(new_n448), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n866), .B2(new_n448), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n448), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT103), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n867), .B1(new_n866), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n866), .A2(new_n882), .A3(new_n448), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n438), .A2(new_n857), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n452), .A2(KEYINPUT104), .B1(new_n434), .B2(new_n443), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n449), .A2(new_n451), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n874), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n876), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n878), .B1(new_n850), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n879), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n843), .B1(new_n901), .B2(new_n674), .ZN(new_n902));
  INV_X1    g0702(.A(new_n900), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n850), .A2(new_n877), .A3(new_n878), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n456), .A3(new_n842), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n456), .B1(new_n729), .B2(new_n732), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n642), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n832), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n731), .B2(new_n831), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(KEYINPUT99), .A3(new_n849), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT99), .ZN(new_n914));
  INV_X1    g0714(.A(new_n831), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n682), .B1(new_n650), .B2(new_n655), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n832), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n849), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n919), .A3(new_n877), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n898), .A2(new_n921), .A3(new_n876), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n875), .B2(new_n876), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n342), .A2(new_n353), .A3(new_n668), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n920), .B1(new_n444), .B2(new_n857), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT105), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n910), .A2(new_n927), .B1(new_n265), .B2(new_n661), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n910), .B2(new_n927), .ZN(new_n929));
  OAI211_X1 g0729(.A(G116), .B(new_n227), .C1(new_n470), .C2(KEYINPUT35), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(KEYINPUT35), .B2(new_n470), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n229), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n276), .A2(G68), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n265), .B(G13), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n929), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NOR2_X1   g0736(.A1(new_n668), .A2(new_n581), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n647), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n602), .B2(new_n937), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT106), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n682), .A2(new_n475), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n512), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n682), .A2(new_n720), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n681), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n945), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n565), .A3(new_n570), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n507), .A2(new_n511), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n682), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n941), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT108), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n948), .A2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(new_n940), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT109), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT109), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n680), .B2(new_n945), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n738), .B(KEYINPUT111), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n945), .A2(new_n683), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT44), .Z(new_n969));
  NOR2_X1   g0769(.A1(new_n945), .A2(new_n683), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n680), .B(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n679), .B1(new_n651), .B2(new_n667), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n681), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n974), .B2(new_n681), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(new_n675), .Z(new_n978));
  AOI22_X1  g0778(.A1(new_n973), .A2(new_n978), .B1(new_n733), .B2(new_n735), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n687), .B(KEYINPUT41), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n967), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n680), .A2(new_n945), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n961), .A2(new_n983), .A3(new_n963), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n965), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n243), .A2(new_n746), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n754), .B1(new_n230), .B2(new_n365), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n798), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n762), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(G68), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n778), .B2(new_n805), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT114), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n287), .B1(new_n201), .B2(new_n776), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G143), .B2(new_n759), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n782), .A2(G159), .B1(new_n765), .B2(G50), .ZN(new_n995));
  INV_X1    g0795(.A(new_n771), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G77), .A2(new_n996), .B1(new_n812), .B2(G137), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n776), .A2(new_n605), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n766), .A2(new_n770), .B1(new_n517), .B2(new_n781), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G107), .C2(new_n989), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n771), .A2(new_n328), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n398), .B(new_n1003), .C1(G317), .C2(new_n812), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT113), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n778), .A2(new_n775), .B1(new_n767), .B2(new_n758), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT112), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1002), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n998), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n756), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n988), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n956), .B2(new_n796), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n985), .A2(new_n1017), .ZN(G387));
  AND2_X1   g0818(.A1(new_n736), .A2(new_n978), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n688), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n736), .B2(new_n978), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n746), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n689), .B(new_n744), .C1(new_n202), .C2(new_n344), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n256), .A2(new_n276), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(KEYINPUT50), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n239), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n744), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n287), .A2(new_n230), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(new_n689), .B1(G107), .B2(new_n230), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT116), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n742), .B1(new_n1035), .B2(new_n754), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n782), .A2(new_n256), .B1(G159), .B2(new_n759), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n276), .B2(new_n778), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n785), .A2(G77), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n398), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n762), .A2(new_n365), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n202), .B2(new_n766), .C1(new_n328), .C2(new_n771), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1038), .B(new_n1043), .C1(G150), .C2(new_n812), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n409), .B1(new_n771), .B2(new_n605), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n759), .A2(G322), .B1(new_n777), .B2(G317), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n767), .B2(new_n781), .C1(new_n775), .C2(new_n766), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT48), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n762), .A2(new_n770), .B1(new_n517), .B2(new_n776), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1045), .B(new_n1051), .C1(G326), .C2(new_n812), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1044), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1036), .B1(new_n1054), .B2(new_n756), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n679), .B2(new_n752), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n978), .B2(new_n966), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1021), .A2(new_n1057), .ZN(G393));
  AOI21_X1  g0858(.A(new_n688), .B1(new_n1019), .B2(new_n973), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n973), .B2(new_n1019), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n973), .A2(new_n966), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n250), .A2(new_n1022), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n753), .B(new_n752), .C1(G97), .C2(new_n686), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n742), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n398), .B1(new_n776), .B2(new_n202), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G77), .B2(new_n989), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n276), .B2(new_n781), .C1(new_n766), .C2(new_n363), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n819), .B(new_n1067), .C1(G143), .C2(new_n812), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n778), .A2(new_n403), .B1(new_n805), .B2(new_n758), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n759), .A2(G317), .B1(new_n777), .B2(G311), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  OAI22_X1  g0872(.A1(new_n766), .A2(new_n517), .B1(new_n775), .B2(new_n781), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n296), .B1(new_n770), .B2(new_n776), .C1(new_n605), .C2(new_n762), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n208), .A2(new_n771), .B1(new_n772), .B2(new_n779), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1068), .A2(new_n1070), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1064), .B1(new_n756), .B2(new_n1077), .C1(new_n949), .C2(new_n796), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1060), .A2(new_n1061), .A3(new_n1078), .ZN(G390));
  NAND2_X1  g0879(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n898), .A2(new_n921), .A3(new_n876), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n925), .B1(new_n917), .B2(new_n918), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n911), .B1(new_n728), .B2(new_n831), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n849), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n925), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n898), .B2(new_n876), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n710), .A2(KEYINPUT89), .A3(G330), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT89), .B1(new_n710), .B2(G330), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n833), .B(new_n849), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1083), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n924), .A2(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n842), .A2(G330), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n849), .A2(new_n833), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1084), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n842), .A2(new_n833), .A3(G330), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n918), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1091), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n833), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1096), .B1(new_n1103), .B2(new_n918), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n917), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n908), .A2(new_n843), .A3(new_n642), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n688), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1098), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1083), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1097), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n908), .A2(new_n843), .A3(new_n642), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n849), .B1(new_n715), .B2(new_n833), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n912), .B1(new_n1115), .B2(new_n1096), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1116), .B2(new_n1102), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT117), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n742), .B1(new_n363), .B2(new_n826), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT118), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  AOI22_X1  g0922(.A1(new_n782), .A2(G137), .B1(new_n765), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  INV_X1    g0924(.A(G132), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n758), .C1(new_n1125), .C2(new_n778), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n776), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT53), .B1(new_n776), .B2(new_n805), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n403), .B2(new_n762), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n287), .B1(new_n771), .B2(new_n276), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G125), .B2(new_n812), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT119), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n296), .B1(new_n416), .B2(new_n776), .C1(new_n766), .C2(new_n328), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n781), .A2(new_n208), .B1(new_n758), .B2(new_n770), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n772), .A2(new_n517), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1134), .A2(new_n811), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n778), .A2(new_n605), .B1(new_n344), .B2(new_n762), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT120), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1130), .A2(new_n1133), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1121), .B1(new_n756), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n924), .B2(new_n750), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1113), .B2(new_n966), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(G378));
  OAI21_X1  g0944(.A(new_n1106), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n317), .A2(new_n665), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n325), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n325), .A2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1147), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1152), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n1150), .A3(new_n1146), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n905), .B2(G330), .ZN(new_n1157));
  OAI211_X1 g0957(.A(G330), .B(new_n1156), .C1(new_n879), .C2(new_n900), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1157), .A2(new_n1159), .A3(new_n926), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1156), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n901), .B2(new_n674), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n444), .A2(new_n857), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n1086), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1162), .A2(new_n1158), .B1(new_n920), .B2(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1145), .A2(KEYINPUT57), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1109), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1112), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1117), .A2(KEYINPUT117), .A3(new_n1092), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1114), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1168), .A2(new_n1175), .A3(new_n687), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1161), .A2(new_n750), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n798), .B1(G50), .B2(new_n827), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n765), .A2(new_n599), .B1(G107), .B2(new_n777), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n605), .B2(new_n758), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n782), .A2(G97), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n398), .A2(G41), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(new_n990), .A3(new_n1039), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n772), .A2(new_n770), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n771), .A2(new_n201), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1180), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT58), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1182), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n276), .C1(G33), .C2(G41), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n759), .A2(G125), .B1(new_n777), .B2(G128), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n804), .B2(new_n766), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n989), .A2(G150), .B1(new_n785), .B2(new_n1122), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1125), .B2(new_n781), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n996), .A2(G159), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n812), .C2(G124), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1190), .B1(KEYINPUT58), .B2(new_n1186), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1178), .B1(new_n1202), .B2(new_n753), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1177), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1174), .B2(new_n967), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1176), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(G375));
  INV_X1    g1011(.A(new_n1105), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n849), .A2(G13), .A3(G33), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n772), .A2(new_n1124), .B1(new_n403), .B2(new_n776), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT123), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n398), .B1(new_n276), .B2(new_n762), .C1(new_n766), .C2(new_n805), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1215), .A2(new_n1185), .A3(new_n1216), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT124), .Z(new_n1218));
  NAND2_X1  g1018(.A1(new_n782), .A2(new_n1122), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n759), .A2(KEYINPUT122), .A3(G132), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n758), .B2(new_n1125), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n777), .A2(G137), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n759), .A2(G294), .B1(new_n777), .B2(G283), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n605), .B2(new_n781), .C1(new_n208), .C2(new_n766), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n287), .B(new_n1041), .C1(G97), .C2(new_n785), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n344), .B2(new_n771), .C1(new_n775), .C2(new_n772), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1218), .A2(new_n1224), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n753), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1230), .B(new_n798), .C1(G68), .C2(new_n827), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1212), .A2(new_n967), .B1(new_n1213), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1116), .A2(new_n1114), .A3(new_n1102), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1107), .A2(new_n1234), .A3(new_n980), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(G381));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1209), .A2(new_n1237), .A3(new_n1210), .ZN(new_n1238));
  INV_X1    g1038(.A(G390), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n839), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G387), .A2(new_n1238), .A3(G381), .A4(new_n1241), .ZN(G407));
  AND3_X1   g1042(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT121), .B1(new_n1176), .B2(new_n1206), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1243), .A2(new_n1244), .A3(G378), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n666), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G407), .A2(G213), .A3(new_n1246), .ZN(G409));
  NAND2_X1  g1047(.A1(new_n1207), .A2(G378), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1107), .A2(new_n687), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1234), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT125), .B1(new_n1234), .B2(new_n1250), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1212), .A2(new_n1253), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1256), .B2(new_n1233), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n839), .B(new_n1232), .C1(new_n1251), .C2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G378), .A2(new_n1205), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1145), .A2(new_n980), .A3(new_n1167), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1260), .A2(new_n1261), .B1(G213), .B2(new_n666), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1248), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1248), .A2(new_n1262), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1259), .B2(KEYINPUT126), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1257), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1258), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1266), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1271), .B(new_n1272), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1265), .A2(new_n1267), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1248), .A2(new_n1277), .A3(new_n1259), .A4(new_n1262), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1264), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1239), .A2(G387), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G390), .A2(new_n1017), .A3(new_n985), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AND2_X1   g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1240), .B2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1240), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1267), .A2(new_n1273), .A3(new_n1270), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1265), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1263), .A2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1282), .B(new_n1285), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1263), .A2(new_n1291), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(G405));
  XNOR2_X1  g1096(.A(new_n1259), .B(KEYINPUT127), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1238), .A2(new_n1248), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1238), .B2(new_n1248), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1287), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1297), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1248), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1245), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1238), .A2(new_n1248), .A3(new_n1297), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1293), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1300), .A2(new_n1305), .ZN(G402));
endmodule


