//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g031(.A1(G113), .A2(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT68), .B1(new_n458), .B2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n459), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n458), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND3_X1  g048(.A1(new_n467), .A2(G2105), .A3(new_n469), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n468), .A2(G112), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n478), .B1(new_n483), .B2(G136), .ZN(G162));
  NAND4_X1  g059(.A1(new_n467), .A2(G138), .A3(new_n468), .A4(new_n469), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AND4_X1   g064(.A1(new_n487), .A2(new_n489), .A3(new_n459), .A4(new_n461), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(KEYINPUT70), .B(G114), .Z(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n468), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n502), .A2(new_n504), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n502), .A2(new_n504), .A3(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(G88), .B1(new_n511), .B2(G50), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n508), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n512), .A2(new_n515), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n513), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n528), .B1(new_n510), .B2(G89), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G51), .A3(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(KEYINPUT7), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT7), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n529), .A2(new_n531), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND3_X1  g115(.A1(new_n530), .A2(new_n513), .A3(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n530), .A2(G52), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n506), .A2(new_n508), .A3(G64), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n501), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n501), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n530), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n509), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n517), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n530), .A2(new_n513), .A3(G91), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n502), .A2(new_n504), .A3(G53), .A4(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n530), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n565), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(G299));
  AOI22_X1  g146(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n542), .B(new_n541), .C1(new_n572), .C2(new_n501), .ZN(G301));
  OAI21_X1  g148(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n530), .A2(G49), .A3(G543), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n509), .ZN(G288));
  NAND3_X1  g152(.A1(new_n530), .A2(G48), .A3(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n511), .A2(new_n580), .A3(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n517), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n510), .A2(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(G305));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  INV_X1    g164(.A(G72), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n517), .A2(new_n589), .B1(new_n590), .B2(new_n505), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n593), .B1(new_n590), .B2(new_n505), .C1(new_n517), .C2(new_n589), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(G651), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n510), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n506), .A2(new_n508), .A3(G66), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(G651), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n511), .A2(G54), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n509), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n530), .A2(new_n513), .A3(KEYINPUT10), .A4(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n609), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n602), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n602), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n566), .B1(new_n621), .B2(new_n501), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n569), .A2(new_n570), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(G868), .B2(new_n624), .ZN(G297));
  OAI21_X1  g200(.A(new_n620), .B1(G868), .B2(new_n624), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n617), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n617), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g207(.A1(new_n468), .A2(G111), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT79), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n467), .A2(G123), .A3(G2105), .A4(new_n469), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(G135), .B2(new_n483), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT15), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2435), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  OAI211_X1 g238(.A(KEYINPUT17), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n662), .ZN(new_n665));
  INV_X1    g240(.A(new_n663), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  OAI221_X1 g243(.A(new_n664), .B1(new_n665), .B2(new_n666), .C1(new_n668), .C2(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n661), .A3(new_n663), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT81), .Z(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(G229));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  NAND3_X1  g274(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n700));
  INV_X1    g275(.A(G129), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n700), .C1(new_n474), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n483), .B2(G141), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G29), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT29), .Z(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G5), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G171), .B2(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G1961), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT95), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G28), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n638), .A2(G29), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G21), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G168), .B2(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G11), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n720), .A2(new_n721), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n723), .A2(G1966), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n708), .B(new_n714), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n554), .B2(new_n734), .ZN(new_n736));
  MUX2_X1   g311(.A(new_n735), .B(new_n736), .S(KEYINPUT88), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G4), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n617), .B2(new_n734), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n716), .A2(G1961), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n737), .B2(G1341), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n734), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n624), .B2(new_n734), .ZN(new_n748));
  INV_X1    g323(.A(G1956), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n742), .A2(new_n744), .A3(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n738), .B(new_n751), .C1(new_n713), .C2(new_n712), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n706), .A2(new_n707), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n459), .A2(new_n461), .A3(G127), .ZN(new_n754));
  NAND2_X1  g329(.A1(G115), .A2(G2104), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n468), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT25), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n483), .B2(G139), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n481), .B2(new_n482), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT90), .B1(new_n763), .B2(new_n758), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n756), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G33), .ZN(new_n767));
  INV_X1    g342(.A(G2072), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n733), .A2(new_n752), .A3(new_n753), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n734), .A2(G24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n600), .B2(new_n734), .ZN(new_n773));
  INV_X1    g348(.A(G1986), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G25), .A2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G119), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n468), .A2(G107), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n474), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n483), .B2(G131), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n776), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G1991), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT83), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n782), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n734), .A2(G6), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n734), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(new_n694), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT84), .B(KEYINPUT32), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT85), .ZN(new_n794));
  XNOR2_X1  g369(.A(G288), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n793), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT86), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n734), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n734), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1971), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n800), .A2(KEYINPUT34), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT34), .B1(new_n800), .B2(new_n804), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n775), .B(new_n786), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT36), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n709), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n709), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT28), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n483), .A2(G140), .ZN(new_n814));
  INV_X1    g389(.A(G128), .ZN(new_n815));
  NOR2_X1   g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT89), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n474), .A2(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n709), .A2(G26), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n813), .B2(new_n823), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2067), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n771), .A2(new_n808), .A3(new_n812), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n767), .A2(new_n768), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT91), .Z(new_n829));
  AND2_X1   g404(.A1(KEYINPUT24), .A2(G34), .ZN(new_n830));
  NOR2_X1   g405(.A1(KEYINPUT24), .A2(G34), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n830), .A2(new_n831), .A3(G29), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n472), .B2(G29), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G2084), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n827), .A2(new_n829), .A3(new_n835), .ZN(G311));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n807), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n826), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(new_n770), .ZN(new_n840));
  INV_X1    g415(.A(new_n829), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n840), .A2(new_n841), .A3(new_n834), .A4(new_n812), .ZN(G150));
  NAND2_X1  g417(.A1(new_n511), .A2(G55), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n530), .A2(new_n513), .A3(G93), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n501), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT98), .B(G860), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n617), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n554), .A2(new_n846), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n511), .A2(G43), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n530), .A2(new_n513), .A3(G81), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n853), .B(new_n854), .C1(new_n548), .C2(new_n501), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n843), .A2(new_n844), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n845), .A2(new_n501), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT39), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n851), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n849), .B1(new_n861), .B2(new_n847), .ZN(G145));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  INV_X1    g438(.A(new_n704), .ZN(new_n864));
  INV_X1    g439(.A(new_n756), .ZN(new_n865));
  INV_X1    g440(.A(new_n764), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n763), .A2(KEYINPUT90), .A3(new_n758), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n499), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n765), .A2(G164), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n869), .A2(new_n821), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n821), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n820), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n869), .A2(new_n821), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n704), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G130), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n468), .A2(G118), .ZN(new_n880));
  OAI22_X1  g455(.A1(new_n474), .A2(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n483), .B2(G142), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n641), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n781), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n873), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n873), .B2(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n863), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(KEYINPUT99), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n472), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(new_n638), .Z(new_n890));
  NAND3_X1  g465(.A1(new_n873), .A2(new_n877), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT100), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  INV_X1    g469(.A(new_n890), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n885), .B2(new_n886), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g473(.A(new_n859), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n629), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n616), .A2(G299), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n624), .A2(new_n610), .A3(new_n609), .A4(new_n615), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT101), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n905), .B1(new_n913), .B2(new_n900), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G303), .B(G305), .ZN(new_n917));
  XNOR2_X1  g492(.A(G288), .B(KEYINPUT85), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n598), .B2(new_n599), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n595), .A2(new_n597), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT77), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n795), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n917), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n917), .B1(new_n923), .B2(new_n919), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n916), .B(new_n926), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n846), .B(new_n927), .S(G868), .Z(G295));
  MUX2_X1   g503(.A(new_n846), .B(new_n927), .S(G868), .Z(G331));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n529), .A2(G301), .A3(new_n531), .A4(new_n538), .ZN(new_n931));
  INV_X1    g506(.A(new_n538), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n530), .A2(new_n513), .A3(G89), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n527), .B1(new_n513), .B2(new_n524), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n527), .A2(new_n506), .A3(new_n508), .A4(new_n524), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n531), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G171), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n899), .A2(new_n930), .A3(new_n931), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n937), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n859), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n852), .A2(new_n931), .A3(new_n937), .A4(new_n858), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(KEYINPUT104), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n910), .A2(new_n912), .A3(new_n938), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n904), .A2(new_n940), .A3(new_n941), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n926), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n926), .A3(new_n947), .A4(new_n944), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n946), .A2(new_n894), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n943), .A2(new_n944), .ZN(new_n953));
  INV_X1    g528(.A(new_n926), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n949), .A2(new_n950), .A3(new_n952), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n940), .A2(new_n941), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n908), .B1(new_n901), .B2(new_n902), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n911), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n942), .A2(new_n938), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n904), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n958), .B(new_n964), .C1(new_n911), .C2(new_n959), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n954), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n946), .A2(new_n967), .A3(new_n894), .A4(new_n948), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n968), .B2(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n946), .A2(new_n955), .A3(new_n894), .A4(new_n948), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT107), .B1(new_n970), .B2(new_n951), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n956), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n956), .A2(new_n969), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n970), .A2(new_n951), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n968), .A2(new_n951), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n957), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT109), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n976), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n490), .B1(new_n485), .B2(KEYINPUT4), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n496), .A2(new_n497), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n465), .A2(G40), .A3(new_n470), .A4(new_n471), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n821), .A2(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n821), .A2(G2067), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n995), .B2(new_n864), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT125), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  INV_X1    g577(.A(new_n992), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n864), .A2(G1996), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n992), .B1(new_n995), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n704), .A2(new_n997), .A3(new_n1003), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1003), .B1(new_n1011), .B2(new_n993), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n781), .A2(new_n785), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1003), .B1(new_n1013), .B2(new_n1010), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n600), .A2(new_n774), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n1003), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1002), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n694), .B1(new_n586), .B2(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n582), .A2(new_n1023), .A3(new_n586), .A4(new_n587), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n991), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n499), .A2(new_n1026), .A3(new_n985), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n918), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT112), .B(G8), .C1(new_n988), .C2(new_n991), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1027), .A2(G8), .A3(new_n1031), .A4(G288), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1036), .B2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1035), .B(new_n1038), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1030), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT45), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n990), .A2(new_n1026), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n991), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n499), .A2(KEYINPUT111), .A3(new_n1046), .A4(new_n985), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1051), .B2(G2090), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G303), .A2(G8), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n1053), .B(KEYINPUT55), .Z(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(G8), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1040), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1026), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1048), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT115), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1065), .A3(new_n1048), .A4(new_n1062), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n713), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1057), .B1(new_n1067), .B2(new_n1044), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1056), .B1(new_n1068), .B2(new_n1054), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1042), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1045), .A2(new_n1047), .A3(new_n1074), .A4(new_n1050), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1042), .A2(new_n1076), .A3(new_n1071), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(G168), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1070), .B1(new_n1078), .B2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1070), .B1(new_n1082), .B2(G286), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1069), .B1(KEYINPUT62), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1051), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n990), .A2(new_n811), .A3(new_n1026), .A4(new_n1041), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n991), .B1(new_n988), .B2(new_n989), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1091), .A2(KEYINPUT53), .A3(new_n811), .A4(new_n1041), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1080), .B(new_n1099), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1085), .A2(KEYINPUT123), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1040), .A2(new_n1055), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1066), .A2(new_n713), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT114), .B1(new_n1058), .B2(new_n1026), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1060), .B(new_n991), .C1(new_n988), .C2(KEYINPUT50), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1065), .B1(new_n1106), .B2(new_n1048), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1044), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1054), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1041), .A2(KEYINPUT53), .A3(new_n811), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1091), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1114), .B2(new_n1091), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(G301), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1111), .A2(new_n1120), .A3(new_n1084), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G299), .B(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1042), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1048), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1104), .A2(new_n1105), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1123), .B(new_n1126), .C1(new_n1128), .C2(G1956), .ZN(new_n1129));
  NOR2_X1   g704(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1123), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1956), .B1(new_n1106), .B2(new_n1048), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1126), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1063), .A2(new_n749), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1027), .A2(G2067), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1051), .B2(new_n741), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1139), .B(new_n616), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n616), .A2(new_n1139), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n617), .A2(KEYINPUT120), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1123), .B1(new_n1136), .B2(new_n1126), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1130), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1027), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1027), .A2(KEYINPUT118), .A3(new_n1152), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1155), .B(new_n1156), .C1(G1996), .C2(new_n1042), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1157), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT59), .B1(new_n1157), .B2(new_n554), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1138), .A2(new_n1149), .A3(new_n1151), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1141), .A2(new_n616), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1129), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT117), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1129), .C1(new_n1150), .C2(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(G171), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1169), .B(KEYINPUT54), .C1(G171), .C2(new_n1093), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1121), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1030), .A2(G1976), .A3(G288), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n694), .B2(new_n788), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1040), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1173), .A2(new_n1028), .B1(new_n1174), .B2(new_n1055), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1082), .A2(G8), .A3(G168), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1069), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1054), .B1(new_n1052), .B2(G8), .ZN(new_n1179));
  OR4_X1    g754(.A1(new_n1176), .A2(new_n1102), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1175), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1083), .A2(new_n1081), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT62), .B1(new_n1182), .B2(new_n1079), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1183), .A2(new_n1100), .A3(new_n1111), .A4(new_n1098), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1101), .A2(new_n1171), .A3(new_n1181), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(G290), .A2(G1986), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1003), .B1(new_n1188), .B2(new_n1016), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1015), .A2(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1187), .A2(KEYINPUT124), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT124), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1020), .B1(new_n1191), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(new_n977), .A2(new_n978), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n676), .A2(G319), .ZN(new_n1196));
  INV_X1    g770(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g773(.A1(G401), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  AOI21_X1  g775(.A(G229), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1202));
  NAND4_X1  g776(.A1(new_n1200), .A2(new_n1201), .A3(new_n897), .A4(new_n1202), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1204));
  NAND4_X1  g778(.A1(new_n897), .A2(new_n659), .A3(new_n1204), .A4(new_n1202), .ZN(G225));
  NAND2_X1  g779(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1206), .ZN(G308));
endmodule


