//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT86), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT87), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(KEYINPUT2), .B2(G113), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n194), .A2(new_n196), .B1(KEYINPUT2), .B2(G113), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n197), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT4), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(KEYINPUT77), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G104), .ZN(new_n209));
  OR2_X1    g023(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(G107), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n200), .B1(new_n201), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT79), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT78), .A2(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT78), .A2(G101), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n204), .B1(new_n206), .B2(new_n205), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT77), .B1(new_n209), .B2(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n220), .B(new_n223), .C1(new_n226), .C2(new_n207), .ZN(new_n227));
  INV_X1    g041(.A(new_n223), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT79), .B1(new_n216), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n226), .B2(new_n207), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT4), .B1(new_n232), .B2(new_n202), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n219), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n216), .A2(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n220), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(KEYINPUT79), .A3(new_n228), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n198), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n239), .A2(G116), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(G113), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT82), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n197), .A2(new_n198), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n248), .A3(G113), .A4(new_n244), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G101), .B1(new_n231), .B2(new_n204), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G122), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n234), .A2(new_n252), .A3(new_n254), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(KEYINPUT6), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT0), .A4(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(G146), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G125), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT1), .B1(new_n261), .B2(G146), .ZN(new_n271));
  OAI211_X1 g085(.A(G128), .B(new_n271), .C1(new_n264), .C2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n260), .B(new_n262), .C1(KEYINPUT1), .C2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G224), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT83), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n253), .A2(new_n283), .A3(new_n255), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n258), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(G113), .A3(new_n244), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n247), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(new_n251), .C1(new_n227), .C2(new_n229), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n254), .B(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n238), .B2(new_n251), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n277), .B(new_n270), .C1(new_n296), .C2(new_n280), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT7), .B1(new_n279), .B2(G953), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n251), .B1(new_n227), .B2(new_n229), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n250), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT84), .A3(new_n290), .A4(new_n291), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n299), .A3(new_n257), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n191), .B1(new_n285), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n303), .A2(new_n304), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n258), .A2(new_n282), .A3(new_n284), .ZN(new_n308));
  INV_X1    g122(.A(new_n190), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G475), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n276), .B2(KEYINPUT71), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(G125), .A3(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(G146), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT72), .B1(new_n318), .B2(new_n259), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n276), .A2(G140), .ZN(new_n321));
  AND4_X1   g135(.A1(KEYINPUT72), .A2(new_n320), .A3(new_n321), .A4(new_n259), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n317), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(KEYINPUT88), .A2(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(KEYINPUT88), .A2(G143), .ZN(new_n325));
  NOR2_X1   g139(.A1(G237), .A2(G953), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n324), .A2(new_n325), .B1(new_n326), .B2(G214), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  INV_X1    g142(.A(G953), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G214), .ZN(new_n330));
  NOR2_X1   g144(.A1(KEYINPUT88), .A2(G143), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT18), .B(G131), .C1(new_n327), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n325), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(new_n331), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(G214), .A3(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n323), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n316), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n320), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n340), .A2(new_n259), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n259), .B1(new_n340), .B2(new_n342), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G131), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n335), .B2(new_n336), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT17), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n327), .A2(new_n332), .A3(G131), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(new_n347), .A3(KEYINPUT17), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n339), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(G113), .B(G122), .Z(new_n353));
  XOR2_X1   g167(.A(KEYINPUT89), .B(G104), .Z(new_n354));
  XOR2_X1   g168(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n355), .B(new_n339), .C1(new_n349), .C2(new_n351), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n312), .B1(new_n359), .B2(new_n304), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n340), .A2(new_n342), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G146), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT19), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n318), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n314), .A2(KEYINPUT19), .A3(new_n316), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n259), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n363), .B(new_n367), .C1(new_n350), .C2(new_n347), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n339), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT90), .A3(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n358), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT90), .B1(new_n369), .B2(new_n356), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT91), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n356), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT90), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n358), .A4(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT20), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n358), .A3(new_n370), .ZN(new_n382));
  NOR3_X1   g196(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(G234), .A2(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(G902), .A3(G953), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT97), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT21), .B(G898), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n329), .A2(G952), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(G234), .B2(G237), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n261), .B2(G128), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n273), .A2(KEYINPUT93), .A3(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n261), .A2(G128), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n395), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n401), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G134), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT94), .A3(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(G116), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT92), .A2(G122), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(G116), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n208), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n413), .ZN(new_n417));
  NOR2_X1   g231(.A1(KEYINPUT92), .A2(G122), .ZN(new_n418));
  OAI21_X1  g232(.A(G116), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n415), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G107), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(KEYINPUT14), .A3(G107), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n419), .A2(KEYINPUT14), .A3(G107), .A4(new_n420), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n405), .A2(new_n408), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT13), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n400), .B1(new_n399), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(new_n406), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n406), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n416), .A3(new_n421), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT9), .B(G234), .ZN(new_n432));
  INV_X1    g246(.A(G217), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n432), .A2(new_n433), .A3(G953), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT95), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT96), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT96), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n425), .A2(new_n430), .A3(new_n436), .A4(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n304), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  AND4_X1   g260(.A1(new_n361), .A2(new_n385), .A3(new_n394), .A4(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G221), .B1(new_n432), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n238), .A2(KEYINPUT10), .A3(new_n275), .A4(new_n251), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n275), .B(new_n251), .C1(new_n227), .C2(new_n229), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT10), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n268), .B1(new_n218), .B2(new_n201), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n230), .B2(new_n233), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT64), .B1(new_n400), .B2(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT11), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT64), .B(new_n458), .C1(new_n400), .C2(G137), .ZN(new_n459));
  INV_X1    g273(.A(G137), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G131), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n456), .B2(KEYINPUT11), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n346), .A3(new_n459), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT80), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n450), .A2(new_n453), .A3(new_n455), .A4(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n329), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n275), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n300), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n451), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT12), .A3(new_n467), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n275), .B1(new_n238), .B2(new_n251), .ZN(new_n479));
  INV_X1    g293(.A(new_n451), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n467), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n474), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n450), .A2(new_n453), .A3(new_n455), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n467), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n473), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n449), .B(new_n304), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n469), .A3(new_n473), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n450), .A2(new_n453), .A3(new_n455), .A4(new_n468), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n483), .B2(new_n478), .ZN(new_n491));
  OAI211_X1 g305(.A(G469), .B(new_n489), .C1(new_n491), .C2(new_n473), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n449), .A2(new_n304), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n311), .A2(new_n447), .A3(new_n448), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n433), .B1(G234), .B2(new_n304), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT74), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n243), .A2(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n273), .A2(G119), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT24), .B(G110), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT23), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n243), .B2(G128), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n273), .A2(KEYINPUT23), .A3(G119), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n500), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n503), .A2(new_n505), .B1(new_n509), .B2(G110), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n320), .A2(new_n321), .A3(new_n259), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n318), .A2(KEYINPUT72), .A3(new_n259), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n363), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n503), .A2(new_n505), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n343), .B2(new_n344), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n509), .A2(KEYINPUT70), .A3(G110), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT70), .B1(new_n509), .B2(G110), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n329), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(KEYINPUT73), .B(new_n516), .C1(new_n518), .C2(new_n521), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n525), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n499), .B1(new_n533), .B2(G902), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n498), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n499), .B(KEYINPUT25), .C1(new_n533), .C2(G902), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n533), .B(KEYINPUT75), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n497), .A2(G902), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n326), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n546));
  XNOR2_X1  g360(.A(new_n197), .B(new_n198), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n268), .B1(new_n464), .B2(new_n466), .ZN(new_n548));
  AND4_X1   g362(.A1(new_n346), .A2(new_n457), .A3(new_n459), .A4(new_n462), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n400), .A2(G137), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n550), .B2(new_n461), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n272), .A2(new_n274), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n346), .B1(new_n465), .B2(new_n459), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n269), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n275), .A2(new_n466), .A3(new_n551), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n200), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n546), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n548), .A2(new_n553), .A3(new_n547), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n545), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT30), .B1(new_n548), .B2(new_n553), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n200), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n558), .A2(new_n544), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT31), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT66), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n570), .B2(new_n547), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR4_X1   g387(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT66), .A4(KEYINPUT31), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n562), .B(new_n568), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT68), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n580));
  INV_X1    g394(.A(new_n576), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n548), .A2(new_n553), .A3(KEYINPUT30), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n564), .B1(new_n556), .B2(new_n557), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n547), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n567), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n572), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT66), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n571), .A2(new_n569), .A3(new_n572), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n562), .A2(new_n568), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n581), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n580), .B1(new_n591), .B2(KEYINPUT32), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n579), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT69), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n562), .A2(new_n568), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n588), .B2(new_n587), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n581), .A2(new_n578), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n575), .A2(KEYINPUT69), .A3(new_n597), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n545), .B1(new_n566), .B2(new_n560), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n559), .A2(new_n561), .A3(new_n545), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT29), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n554), .A2(new_n558), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n561), .B1(KEYINPUT28), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT29), .A3(new_n544), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n304), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n600), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n540), .B1(new_n593), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n496), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n221), .A2(new_n222), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n612), .B(new_n613), .Z(G3));
  AND2_X1   g428(.A1(new_n495), .A2(new_n448), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n596), .B2(G902), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n577), .A3(new_n540), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n309), .B1(new_n307), .B2(new_n308), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n187), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n438), .B1(new_n431), .B2(KEYINPUT98), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n623), .B(new_n435), .C1(new_n425), .C2(new_n430), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT33), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n440), .A2(new_n626), .A3(new_n441), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n625), .A2(G478), .A3(new_n304), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n442), .A2(new_n443), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n380), .A2(KEYINPUT20), .B1(new_n382), .B2(new_n383), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n630), .B(new_n394), .C1(new_n631), .C2(new_n360), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n618), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n190), .B1(new_n285), .B2(new_n305), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n188), .B1(new_n634), .B2(new_n310), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n630), .B1(new_n631), .B2(new_n360), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n635), .A2(KEYINPUT99), .A3(new_n394), .A4(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n617), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT20), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n373), .A2(new_n379), .A3(new_n644), .A4(new_n374), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n381), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n373), .A2(new_n379), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(KEYINPUT101), .A3(new_n644), .A4(new_n374), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n442), .A2(new_n444), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n442), .A2(new_n444), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n360), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n646), .A2(new_n649), .A3(new_n394), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n635), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n617), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  OAI221_X1 g474(.A(new_n517), .B1(new_n519), .B2(new_n520), .C1(new_n343), .C2(new_n344), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT73), .B1(new_n661), .B2(new_n516), .ZN(new_n662));
  INV_X1    g476(.A(new_n530), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n532), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n664), .B2(new_n526), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n535), .B1(new_n665), .B2(KEYINPUT74), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n497), .A3(new_n537), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n531), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n539), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n673));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n577), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n615), .A2(new_n676), .A3(new_n447), .A4(new_n311), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  OAI211_X1 g493(.A(new_n635), .B(new_n671), .C1(new_n593), .C2(new_n610), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n392), .B(KEYINPUT104), .Z(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n388), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n495), .A3(new_n448), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n273), .ZN(G30));
  NAND2_X1  g502(.A1(new_n306), .A2(new_n310), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT38), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(KEYINPUT38), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n631), .A2(new_n360), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n446), .A4(new_n188), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n685), .B(KEYINPUT39), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n615), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n566), .A2(new_n560), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n545), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n304), .B1(new_n605), .B2(new_n544), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n599), .A3(new_n600), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n672), .B1(new_n704), .B2(new_n593), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n697), .A3(new_n698), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  OAI211_X1 g522(.A(new_n671), .B(new_n187), .C1(new_n619), .C2(new_n620), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n579), .A2(new_n592), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n599), .A2(new_n600), .A3(new_n609), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n630), .B(new_n685), .C1(new_n631), .C2(new_n360), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n448), .A3(new_n495), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n486), .A2(new_n469), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n472), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT12), .B1(new_n477), .B2(new_n467), .ZN(new_n721));
  INV_X1    g535(.A(new_n467), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n482), .B(new_n722), .C1(new_n476), .C2(new_n451), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n469), .B(new_n473), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n449), .B1(new_n725), .B2(new_n304), .ZN(new_n726));
  AOI211_X1 g540(.A(G469), .B(G902), .C1(new_n720), .C2(new_n724), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n728), .B2(new_n448), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n483), .A2(new_n478), .ZN(new_n730));
  INV_X1    g544(.A(new_n474), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n730), .A2(new_n731), .B1(new_n719), .B2(new_n472), .ZN(new_n732));
  OAI21_X1  g546(.A(G469), .B1(new_n732), .B2(G902), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n448), .A4(new_n488), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n638), .A2(new_n633), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT75), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n533), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n533), .A2(new_n738), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n539), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n667), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n710), .B2(new_n711), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n736), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NOR2_X1   g560(.A1(new_n656), .A2(new_n654), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n736), .A2(new_n747), .A3(new_n743), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NAND3_X1  g563(.A1(new_n728), .A2(new_n447), .A3(new_n448), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n680), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n243), .ZN(G21));
  NAND2_X1  g566(.A1(new_n634), .A2(new_n310), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n446), .B1(new_n385), .B2(new_n361), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n394), .A3(new_n187), .A4(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n729), .A2(new_n735), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n673), .B2(new_n674), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT108), .B(G472), .C1(new_n596), .C2(G902), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n545), .B1(new_n606), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n606), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n589), .A2(new_n568), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n576), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n540), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n540), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n756), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NAND3_X1  g586(.A1(new_n728), .A2(new_n635), .A3(new_n448), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n760), .A2(new_n714), .A3(new_n671), .A4(new_n765), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n276), .ZN(G27));
  OAI221_X1 g590(.A(new_n609), .B1(new_n596), .B2(new_n598), .C1(KEYINPUT32), .C2(new_n591), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n540), .ZN(new_n778));
  INV_X1    g592(.A(new_n191), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n307), .B2(new_n308), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n448), .A2(new_n187), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n619), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n492), .A2(KEYINPUT110), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n469), .B1(new_n721), .B2(new_n723), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n472), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n786), .A3(G469), .A4(new_n489), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n488), .A3(new_n494), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n778), .A2(new_n789), .A3(new_n790), .A4(new_n713), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n611), .A2(new_n789), .A3(new_n713), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT111), .B1(new_n792), .B2(KEYINPUT42), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n782), .A2(new_n788), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n743), .A2(new_n794), .A3(new_n714), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n790), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n791), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT112), .B(G131), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G33));
  AND2_X1   g614(.A1(new_n681), .A2(new_n685), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n743), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND3_X1  g617(.A1(new_n306), .A2(new_n310), .A3(new_n187), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n693), .A2(new_n630), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n675), .A3(new_n671), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n785), .A2(new_n489), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n449), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n785), .A2(KEYINPUT45), .A3(new_n489), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n493), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(KEYINPUT46), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n488), .B1(new_n816), .B2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n448), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  INV_X1    g634(.A(new_n695), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n819), .B2(new_n821), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n811), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(new_n460), .ZN(G39));
  NAND3_X1  g640(.A1(new_n711), .A2(new_n592), .A3(new_n579), .ZN(new_n827));
  OR4_X1    g641(.A1(new_n827), .A2(new_n540), .A3(new_n713), .A4(new_n804), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n819), .A2(new_n829), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(new_n313), .ZN(G42));
  AND3_X1   g647(.A1(new_n692), .A2(new_n693), .A3(new_n630), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n704), .A2(new_n593), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n742), .A2(new_n781), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT114), .Z(new_n837));
  XNOR2_X1  g651(.A(new_n728), .B(KEYINPUT49), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n685), .A2(new_n448), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n788), .A2(new_n635), .A3(new_n754), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n706), .A2(new_n843), .B1(new_n712), .B2(new_n716), .ZN(new_n844));
  INV_X1    g658(.A(new_n686), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n671), .A2(new_n760), .A3(new_n714), .A4(new_n765), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n733), .A2(new_n448), .A3(new_n488), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n621), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n712), .A2(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n840), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n705), .A2(new_n842), .B1(new_n680), .B2(new_n715), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n680), .A2(new_n686), .B1(new_n773), .B2(new_n774), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT52), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n844), .A2(new_n849), .A3(new_n840), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT52), .B1(new_n851), .B2(new_n852), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n791), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n792), .A2(KEYINPUT111), .A3(KEYINPUT42), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n796), .B1(new_n795), .B2(new_n790), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n751), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n744), .A2(new_n771), .A3(new_n748), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n689), .A2(new_n495), .A3(new_n448), .A4(new_n187), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n636), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n630), .B(KEYINPUT115), .C1(new_n631), .C2(new_n360), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n540), .A2(new_n577), .A3(new_n394), .A4(new_n616), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n866), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT116), .B1(new_n612), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n868), .A2(new_n869), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n675), .A2(new_n742), .A3(new_n393), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n615), .A3(new_n311), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n876), .B(new_n877), .C1(new_n611), .C2(new_n496), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n446), .B(KEYINPUT117), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n879), .A2(new_n693), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n615), .A2(new_n880), .A3(new_n875), .A4(new_n311), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(new_n677), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n873), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n846), .A2(new_n794), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n804), .A2(new_n672), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n646), .A2(new_n649), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n361), .A2(new_n685), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n879), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n827), .A2(new_n885), .A3(new_n888), .A4(new_n615), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n802), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n863), .A2(new_n865), .A3(new_n883), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n859), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n855), .A2(new_n894), .A3(new_n857), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n855), .B2(new_n857), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n847), .A2(new_n898), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n827), .A2(new_n899), .A3(new_n540), .A4(new_n734), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n751), .B1(new_n900), .B2(new_n737), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n890), .A2(new_n901), .A3(new_n748), .A4(new_n771), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n873), .A2(new_n878), .A3(new_n882), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n798), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n897), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n893), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n892), .B1(new_n859), .B2(new_n891), .ZN(new_n907));
  INV_X1    g721(.A(new_n896), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n855), .A2(new_n894), .A3(new_n857), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  INV_X1    g728(.A(new_n807), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n682), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n770), .ZN(new_n917));
  INV_X1    g731(.A(new_n847), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n692), .A2(new_n188), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT50), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n770), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT50), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT121), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n804), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n830), .A2(new_n831), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n726), .A2(new_n727), .A3(new_n448), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n926), .B(new_n917), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n926), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n915), .A2(new_n930), .A3(new_n682), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n760), .A2(new_n671), .A3(new_n765), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n835), .A2(new_n540), .A3(new_n392), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n930), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n631), .A2(new_n630), .A3(new_n360), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n931), .A2(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n929), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n921), .A2(new_n924), .A3(KEYINPUT121), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n914), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n391), .B1(new_n934), .B2(new_n637), .ZN(new_n940));
  INV_X1    g754(.A(new_n778), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT48), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n931), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n931), .B2(new_n941), .ZN(new_n944));
  OAI221_X1 g758(.A(new_n940), .B1(new_n773), .B2(new_n922), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT50), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n923), .B1(new_n922), .B2(new_n919), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n914), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n929), .A2(new_n948), .A3(new_n936), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n929), .A2(new_n948), .A3(KEYINPUT122), .A4(new_n936), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n939), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n913), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(G952), .A2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n839), .B1(new_n954), .B2(new_n955), .ZN(G75));
  NAND2_X1  g770(.A1(new_n258), .A2(new_n284), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n282), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT124), .B(KEYINPUT55), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n304), .B1(new_n907), .B2(new_n910), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n190), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT56), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n329), .A2(G952), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n960), .A2(new_n963), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n961), .B2(new_n191), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(G51));
  XNOR2_X1  g782(.A(new_n493), .B(KEYINPUT57), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n911), .B1(new_n907), .B2(new_n910), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n725), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n961), .A2(new_n815), .A3(new_n814), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(G54));
  NAND2_X1  g789(.A1(KEYINPUT58), .A2(G475), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n961), .A2(new_n648), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n648), .B1(new_n961), .B2(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n965), .ZN(G60));
  AND2_X1   g794(.A1(new_n625), .A2(new_n627), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n982));
  NAND2_X1  g796(.A1(G478), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n981), .B1(new_n913), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n981), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n970), .B2(new_n971), .ZN(new_n987));
  INV_X1    g801(.A(new_n965), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n985), .A2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR4_X1   g807(.A1(new_n891), .A2(new_n895), .A3(new_n892), .A4(new_n896), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT53), .B1(new_n997), .B2(new_n904), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n993), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n538), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(KEYINPUT126), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n992), .B1(new_n907), .B2(new_n910), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n538), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n965), .B1(new_n1003), .B2(new_n669), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .A4(KEYINPUT61), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n669), .B(new_n993), .C1(new_n994), .C2(new_n998), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n988), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1003), .A2(new_n538), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1006), .A2(new_n1011), .ZN(G66));
  OAI21_X1  g826(.A(G953), .B1(new_n389), .B2(new_n279), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n865), .A2(new_n883), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n957), .B1(G898), .B2(new_n329), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G69));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  INV_X1    g832(.A(new_n717), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n852), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n849), .A2(KEYINPUT127), .A3(new_n717), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n825), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n802), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n832), .A2(new_n798), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n823), .A2(new_n824), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1026), .A2(new_n635), .A3(new_n754), .A4(new_n941), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n329), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n365), .A2(new_n366), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n570), .B(new_n1030), .Z(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(G900), .B2(G953), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n329), .B1(G227), .B2(G900), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n874), .A2(new_n880), .ZN(new_n1037));
  NOR4_X1   g851(.A1(new_n1037), .A2(new_n696), .A3(new_n611), .A4(new_n804), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n825), .A2(new_n832), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1022), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT62), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1040), .A2(new_n1041), .A3(new_n707), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n707), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1039), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g859(.A1(new_n1045), .A2(new_n329), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1034), .B(new_n1036), .C1(new_n1046), .C2(new_n1031), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1033), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1048), .B1(new_n1028), .B2(new_n329), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1031), .B1(new_n1045), .B2(new_n329), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1035), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1047), .A2(new_n1051), .ZN(G72));
  NAND2_X1  g866(.A1(new_n699), .A2(new_n545), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1028), .A2(new_n1014), .ZN(new_n1054));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1039), .A2(new_n1044), .A3(new_n1014), .A4(new_n1042), .ZN(new_n1058));
  AOI211_X1 g872(.A(new_n545), .B(new_n699), .C1(new_n1058), .C2(new_n1056), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n893), .A2(new_n905), .ZN(new_n1060));
  OAI21_X1  g874(.A(new_n1056), .B1(new_n602), .B2(new_n571), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n988), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g876(.A1(new_n1057), .A2(new_n1059), .A3(new_n1062), .ZN(G57));
endmodule


