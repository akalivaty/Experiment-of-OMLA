

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U551 ( .A(n713), .Z(n517) );
  AND2_X1 U552 ( .A1(n790), .A2(n789), .ZN(n805) );
  AND2_X1 U553 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U554 ( .A(n739), .B(KEYINPUT97), .ZN(n713) );
  AND2_X1 U555 ( .A1(n687), .A2(n686), .ZN(n764) );
  NAND2_X2 U556 ( .A1(n689), .A2(n765), .ZN(n739) );
  NOR2_X1 U557 ( .A1(n692), .A2(n691), .ZN(n707) );
  NOR2_X1 U558 ( .A1(n707), .A2(n968), .ZN(n694) );
  NOR2_X1 U559 ( .A1(G651), .A2(n622), .ZN(n644) );
  OR2_X1 U560 ( .A1(n568), .A2(n519), .ZN(n518) );
  AND2_X1 U561 ( .A1(n644), .A2(G43), .ZN(n519) );
  XOR2_X1 U562 ( .A(KEYINPUT70), .B(n564), .Z(n520) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n749) );
  INV_X1 U564 ( .A(G2105), .ZN(n526) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n645) );
  OR2_X1 U567 ( .A1(n569), .A2(n518), .ZN(n984) );
  INV_X1 U568 ( .A(KEYINPUT64), .ZN(n525) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n521), .Z(n874) );
  NAND2_X1 U571 ( .A1(G137), .A2(n874), .ZN(n523) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U573 ( .A1(G113), .A2(n879), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U575 ( .A(n525), .B(n524), .ZN(n688) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n526), .ZN(n877) );
  NAND2_X1 U577 ( .A1(n877), .A2(G125), .ZN(n687) );
  AND2_X1 U578 ( .A1(n688), .A2(n687), .ZN(n528) );
  AND2_X1 U579 ( .A1(n526), .A2(G2104), .ZN(n873) );
  NAND2_X1 U580 ( .A1(G101), .A2(n873), .ZN(n527) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n527), .Z(n685) );
  AND2_X1 U582 ( .A1(n528), .A2(n685), .ZN(G160) );
  XOR2_X1 U583 ( .A(G2443), .B(G2446), .Z(n530) );
  XNOR2_X1 U584 ( .A(G2427), .B(G2451), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n530), .B(n529), .ZN(n536) );
  XOR2_X1 U586 ( .A(G2430), .B(G2454), .Z(n532) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n531) );
  XNOR2_X1 U588 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U589 ( .A(G2435), .B(G2438), .Z(n533) );
  XNOR2_X1 U590 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U591 ( .A(n536), .B(n535), .Z(n537) );
  AND2_X1 U592 ( .A1(G14), .A2(n537), .ZN(G401) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G57), .ZN(G237) );
  INV_X1 U595 ( .A(G108), .ZN(G238) );
  INV_X1 U596 ( .A(G82), .ZN(G220) );
  NAND2_X1 U597 ( .A1(G102), .A2(n873), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G138), .A2(n874), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G114), .A2(n879), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G126), .A2(n877), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n543), .A2(n542), .ZN(G164) );
  NAND2_X1 U604 ( .A1(G89), .A2(n645), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT73), .B(n544), .Z(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT4), .ZN(n548) );
  XNOR2_X1 U607 ( .A(G651), .B(KEYINPUT65), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n622), .A2(n550), .ZN(n546) );
  XNOR2_X2 U609 ( .A(KEYINPUT66), .B(n546), .ZN(n652) );
  NAND2_X1 U610 ( .A1(G76), .A2(n652), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U612 ( .A(KEYINPUT5), .B(n549), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G51), .A2(n644), .ZN(n554) );
  XNOR2_X1 U614 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n552) );
  NOR2_X1 U615 ( .A1(G543), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n648) );
  NAND2_X1 U617 ( .A1(G63), .A2(n648), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(KEYINPUT7), .B(n559), .ZN(G168) );
  XNOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n834) );
  NAND2_X1 U628 ( .A1(n834), .A2(G567), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n562), .Z(G234) );
  NAND2_X1 U630 ( .A1(n645), .A2(G81), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n563), .Z(n565) );
  NAND2_X1 U632 ( .A1(n652), .A2(G68), .ZN(n564) );
  NOR2_X1 U633 ( .A1(n565), .A2(n520), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n648), .A2(G56), .ZN(n567) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n567), .Z(n568) );
  XNOR2_X1 U637 ( .A(G860), .B(KEYINPUT71), .ZN(n595) );
  OR2_X1 U638 ( .A1(n984), .A2(n595), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G77), .A2(n652), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G90), .A2(n645), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U642 ( .A(KEYINPUT9), .B(n572), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n648), .A2(G64), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G52), .A2(n644), .ZN(n573) );
  AND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G92), .A2(n645), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G54), .A2(n644), .ZN(n578) );
  NAND2_X1 U650 ( .A1(G66), .A2(n648), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n652), .A2(G79), .ZN(n579) );
  XOR2_X1 U653 ( .A(KEYINPUT72), .B(n579), .Z(n580) );
  NOR2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n584), .B(KEYINPUT15), .ZN(n901) );
  INV_X1 U657 ( .A(n901), .ZN(n979) );
  INV_X1 U658 ( .A(G868), .ZN(n663) );
  NAND2_X1 U659 ( .A1(n979), .A2(n663), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G78), .A2(n652), .ZN(n588) );
  NAND2_X1 U662 ( .A1(G53), .A2(n644), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n645), .A2(G91), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G65), .A2(n648), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n968) );
  INV_X1 U668 ( .A(n968), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G286), .A2(n663), .ZN(n594) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n596), .A2(n901), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n984), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G868), .A2(n901), .ZN(n598) );
  NOR2_X1 U677 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n601), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G99), .A2(n873), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G111), .A2(n879), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U683 ( .A(KEYINPUT78), .B(n604), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G123), .A2(n877), .ZN(n605) );
  XOR2_X1 U685 ( .A(KEYINPUT77), .B(n605), .Z(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U687 ( .A1(G135), .A2(n874), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n923) );
  XNOR2_X1 U690 ( .A(n923), .B(G2096), .ZN(n612) );
  INV_X1 U691 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n645), .A2(G93), .ZN(n614) );
  NAND2_X1 U694 ( .A1(G67), .A2(n648), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G80), .A2(n652), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G55), .A2(n644), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n664) );
  NAND2_X1 U700 ( .A1(G559), .A2(n901), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n984), .B(n619), .ZN(n661) );
  NOR2_X1 U702 ( .A1(G860), .A2(n661), .ZN(n620) );
  XOR2_X1 U703 ( .A(KEYINPUT79), .B(n620), .Z(n621) );
  XOR2_X1 U704 ( .A(n664), .B(n621), .Z(G145) );
  NAND2_X1 U705 ( .A1(G87), .A2(n622), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n648), .A2(n625), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n644), .A2(G49), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G73), .A2(n652), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n628), .B(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G48), .A2(n644), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G61), .A2(n648), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n645), .A2(G86), .ZN(n631) );
  XOR2_X1 U717 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U720 ( .A1(n645), .A2(G88), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G75), .A2(n652), .ZN(n637) );
  NAND2_X1 U722 ( .A1(G62), .A2(n648), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G50), .A2(n644), .ZN(n638) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n638), .ZN(n639) );
  NOR2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U728 ( .A(KEYINPUT82), .B(n643), .Z(G166) );
  NAND2_X1 U729 ( .A1(G47), .A2(n644), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G85), .A2(n645), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n648), .A2(G60), .ZN(n649) );
  XOR2_X1 U733 ( .A(KEYINPUT68), .B(n649), .Z(n650) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n652), .A2(G72), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n654), .A2(n653), .ZN(G290) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n656) );
  XNOR2_X1 U738 ( .A(G288), .B(n968), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n656), .B(n655), .ZN(n658) );
  XOR2_X1 U740 ( .A(G305), .B(G166), .Z(n657) );
  XNOR2_X1 U741 ( .A(n658), .B(n657), .ZN(n660) );
  XOR2_X1 U742 ( .A(G290), .B(n664), .Z(n659) );
  XNOR2_X1 U743 ( .A(n660), .B(n659), .ZN(n904) );
  XNOR2_X1 U744 ( .A(n904), .B(n661), .ZN(n662) );
  NOR2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U746 ( .A1(G868), .A2(n664), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n666), .A2(n665), .ZN(G295) );
  XOR2_X1 U748 ( .A(KEYINPUT21), .B(KEYINPUT84), .Z(n670) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U751 ( .A1(n668), .A2(G2090), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U753 ( .A(KEYINPUT85), .B(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(KEYINPUT86), .B(G44), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n673), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U757 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U759 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n674) );
  XNOR2_X1 U760 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U761 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G96), .A2(n677), .ZN(n838) );
  NAND2_X1 U763 ( .A1(n838), .A2(G2106), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U765 ( .A1(G237), .A2(n678), .ZN(n679) );
  XOR2_X1 U766 ( .A(KEYINPUT88), .B(n679), .Z(n680) );
  NOR2_X1 U767 ( .A1(G238), .A2(n680), .ZN(n681) );
  XNOR2_X1 U768 ( .A(KEYINPUT89), .B(n681), .ZN(n839) );
  NAND2_X1 U769 ( .A1(n839), .A2(G567), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n915) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n915), .A2(n684), .ZN(n837) );
  NAND2_X1 U773 ( .A1(n837), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G301), .ZN(G171) );
  XOR2_X1 U775 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  XNOR2_X1 U776 ( .A(G1981), .B(G305), .ZN(n989) );
  AND2_X1 U777 ( .A1(G40), .A2(n685), .ZN(n686) );
  AND2_X1 U778 ( .A1(n688), .A2(n764), .ZN(n689) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n765) );
  NAND2_X1 U780 ( .A1(n517), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  INV_X1 U782 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U783 ( .A1(n997), .A2(n517), .ZN(n691) );
  XOR2_X1 U784 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n693) );
  XNOR2_X1 U785 ( .A(n694), .B(n693), .ZN(n711) );
  INV_X1 U786 ( .A(G1996), .ZN(n695) );
  NOR2_X1 U787 ( .A1(n739), .A2(n695), .ZN(n696) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U789 ( .A1(n739), .A2(G1341), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n984), .A2(n699), .ZN(n700) );
  OR2_X1 U792 ( .A1(n901), .A2(n700), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n901), .A2(n700), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n517), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n739), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n707), .A2(n968), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U802 ( .A(n712), .B(KEYINPUT29), .ZN(n717) );
  INV_X1 U803 ( .A(G1961), .ZN(n996) );
  NAND2_X1 U804 ( .A1(n996), .A2(n739), .ZN(n715) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U806 ( .A1(n517), .A2(n955), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n719) );
  AND2_X1 U808 ( .A1(G171), .A2(n719), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT99), .ZN(n736) );
  NOR2_X1 U811 ( .A1(G171), .A2(n719), .ZN(n724) );
  NAND2_X1 U812 ( .A1(G8), .A2(n739), .ZN(n798) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n798), .ZN(n727) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n739), .ZN(n728) );
  NOR2_X1 U815 ( .A1(n727), .A2(n728), .ZN(n720) );
  NAND2_X1 U816 ( .A1(G8), .A2(n720), .ZN(n721) );
  XNOR2_X1 U817 ( .A(KEYINPUT30), .B(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(G168), .A2(n722), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n726) );
  XOR2_X1 U820 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n725) );
  XNOR2_X1 U821 ( .A(n726), .B(n725), .ZN(n735) );
  AND2_X1 U822 ( .A1(n736), .A2(n735), .ZN(n733) );
  INV_X1 U823 ( .A(n727), .ZN(n731) );
  NAND2_X1 U824 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n729), .B(KEYINPUT96), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U828 ( .A(n734), .B(KEYINPUT101), .Z(n752) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n738) );
  AND2_X1 U830 ( .A1(G286), .A2(G8), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n748) );
  INV_X1 U832 ( .A(G8), .ZN(n746) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n739), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n740), .B(KEYINPUT102), .ZN(n742) );
  NOR2_X1 U835 ( .A1(n798), .A2(G1971), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U837 ( .A(KEYINPUT103), .B(n743), .Z(n744) );
  NAND2_X1 U838 ( .A1(n744), .A2(G303), .ZN(n745) );
  OR2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U840 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n791) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NOR2_X1 U843 ( .A1(n791), .A2(n976), .ZN(n755) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n753) );
  XOR2_X1 U845 ( .A(KEYINPUT104), .B(n753), .Z(n970) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U847 ( .A1(n970), .A2(n759), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G288), .A2(G1976), .ZN(n756) );
  XOR2_X1 U850 ( .A(KEYINPUT105), .B(n756), .Z(n969) );
  INV_X1 U851 ( .A(n798), .ZN(n757) );
  NAND2_X1 U852 ( .A1(n969), .A2(n757), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n989), .A2(n762), .ZN(n790) );
  NOR2_X1 U856 ( .A1(n798), .A2(n970), .ZN(n763) );
  NAND2_X1 U857 ( .A1(KEYINPUT33), .A2(n763), .ZN(n788) );
  NAND2_X1 U858 ( .A1(n688), .A2(n764), .ZN(n766) );
  NOR2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n829) );
  INV_X1 U860 ( .A(n829), .ZN(n787) );
  XNOR2_X1 U861 ( .A(G1986), .B(G290), .ZN(n972) );
  NAND2_X1 U862 ( .A1(G105), .A2(n873), .ZN(n767) );
  XNOR2_X1 U863 ( .A(n767), .B(KEYINPUT38), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G141), .A2(n874), .ZN(n769) );
  NAND2_X1 U865 ( .A1(G117), .A2(n879), .ZN(n768) );
  NAND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U867 ( .A1(G129), .A2(n877), .ZN(n770) );
  XNOR2_X1 U868 ( .A(KEYINPUT93), .B(n770), .ZN(n771) );
  NOR2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U871 ( .A(KEYINPUT94), .B(n775), .ZN(n886) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n886), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G131), .A2(n874), .ZN(n776) );
  XOR2_X1 U874 ( .A(KEYINPUT92), .B(n776), .Z(n781) );
  NAND2_X1 U875 ( .A1(G107), .A2(n879), .ZN(n778) );
  NAND2_X1 U876 ( .A1(G119), .A2(n877), .ZN(n777) );
  NAND2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U878 ( .A(KEYINPUT91), .B(n779), .Z(n780) );
  NOR2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n873), .A2(G95), .ZN(n782) );
  NAND2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n890) );
  NAND2_X1 U882 ( .A1(G1991), .A2(n890), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n785), .A2(n784), .ZN(n920) );
  NOR2_X1 U884 ( .A1(n972), .A2(n920), .ZN(n786) );
  OR2_X1 U885 ( .A1(n787), .A2(n786), .ZN(n803) );
  AND2_X1 U886 ( .A1(n788), .A2(n803), .ZN(n789) );
  INV_X1 U887 ( .A(n791), .ZN(n794) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U889 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n798), .A2(n795), .ZN(n801) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U893 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  NOR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U895 ( .A(KEYINPUT95), .B(n799), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  AND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X2 U898 ( .A1(n805), .A2(n804), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G104), .A2(n873), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G140), .A2(n874), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n808), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G116), .A2(n879), .ZN(n810) );
  NAND2_X1 U904 ( .A1(G128), .A2(n877), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U908 ( .A(KEYINPUT36), .B(n814), .Z(n898) );
  XOR2_X1 U909 ( .A(G2067), .B(KEYINPUT37), .Z(n817) );
  AND2_X1 U910 ( .A1(n898), .A2(n817), .ZN(n937) );
  NAND2_X1 U911 ( .A1(n829), .A2(n937), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n815), .A2(n824), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n816), .B(KEYINPUT106), .ZN(n832) );
  NOR2_X1 U914 ( .A1(n898), .A2(n817), .ZN(n921) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n886), .ZN(n930) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n890), .ZN(n924) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XOR2_X1 U918 ( .A(n818), .B(KEYINPUT107), .Z(n819) );
  NOR2_X1 U919 ( .A1(n924), .A2(n819), .ZN(n820) );
  XNOR2_X1 U920 ( .A(n820), .B(KEYINPUT108), .ZN(n821) );
  NOR2_X1 U921 ( .A1(n920), .A2(n821), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n930), .A2(n822), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U925 ( .A(KEYINPUT109), .B(n826), .ZN(n827) );
  NOR2_X1 U926 ( .A1(n921), .A2(n827), .ZN(n828) );
  XOR2_X1 U927 ( .A(KEYINPUT110), .B(n828), .Z(n830) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U933 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U935 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n841) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2072), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U945 ( .A(n842), .B(G2100), .Z(n844) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2084), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U949 ( .A(G2678), .B(KEYINPUT111), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U951 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U952 ( .A(G1966), .B(G1971), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1981), .B(G1976), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n851), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U958 ( .A(G2474), .B(G1956), .Z(n855) );
  XNOR2_X1 U959 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G100), .A2(n873), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G112), .A2(n879), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G124), .A2(n877), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n860), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G136), .A2(n874), .ZN(n861) );
  XNOR2_X1 U968 ( .A(n861), .B(KEYINPUT112), .ZN(n862) );
  NAND2_X1 U969 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U970 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G118), .A2(n879), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G130), .A2(n877), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G106), .A2(n873), .ZN(n869) );
  NAND2_X1 U975 ( .A1(G142), .A2(n874), .ZN(n868) );
  NAND2_X1 U976 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  NOR2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G103), .A2(n873), .ZN(n876) );
  NAND2_X1 U980 ( .A1(G139), .A2(n874), .ZN(n875) );
  NAND2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n877), .A2(G127), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n878), .Z(n881) );
  NAND2_X1 U984 ( .A1(n879), .A2(G115), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n916) );
  XOR2_X1 U988 ( .A(n885), .B(n916), .Z(n888) );
  XNOR2_X1 U989 ( .A(G160), .B(n886), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U991 ( .A(n923), .B(G162), .Z(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(n892), .B(n891), .Z(n897) );
  XOR2_X1 U994 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U997 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U1001 ( .A(KEYINPUT116), .B(G286), .Z(n903) );
  XNOR2_X1 U1002 ( .A(G171), .B(n901), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n984), .B(n904), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n915), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT117), .B(n910), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n915), .ZN(G319) );
  XOR2_X1 U1017 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n919), .Z(n940) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n935) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT119), .B(n922), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(KEYINPUT120), .B(n927), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G162), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(KEYINPUT121), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n931), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT122), .B(n938), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n964), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1040 ( .A(KEYINPUT123), .B(G2090), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(G35), .ZN(n962) );
  XNOR2_X1 U1042 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1044 ( .A(G32), .B(G1996), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(n946), .B(KEYINPUT125), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(G28), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G25), .B(G1991), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1054 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n958), .B(KEYINPUT53), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n964), .B(n963), .ZN(n966) );
  INV_X1 U1060 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n967), .ZN(n1023) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(n968), .B(G1956), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n983) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G171), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1348), .B(n979), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(KEYINPUT127), .B(n987), .Z(n993) );
  XOR2_X1 U1078 ( .A(G1966), .B(G168), .Z(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1080 ( .A(KEYINPUT57), .B(n990), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT126), .B(n991), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n1021) );
  INV_X1 U1084 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1085 ( .A(G5), .B(n996), .ZN(n1009) );
  XNOR2_X1 U1086 ( .A(G20), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT59), .B(G1348), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(G1976), .B(G23), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

