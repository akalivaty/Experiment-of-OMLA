

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  XOR2_X1 U322 ( .A(n345), .B(n344), .Z(n290) );
  XOR2_X1 U323 ( .A(n340), .B(n366), .Z(n291) );
  INV_X1 U324 ( .A(KEYINPUT46), .ZN(n391) );
  INV_X1 U325 ( .A(n461), .ZN(n420) );
  XNOR2_X1 U326 ( .A(n395), .B(KEYINPUT113), .ZN(n396) );
  XNOR2_X1 U327 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U328 ( .A(n346), .B(n290), .ZN(n353) );
  XNOR2_X1 U329 ( .A(n353), .B(n352), .ZN(n578) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n456) );
  XNOR2_X1 U331 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT79), .B(KEYINPUT11), .Z(n293) );
  XNOR2_X1 U334 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U336 ( .A(KEYINPUT80), .B(KEYINPUT65), .Z(n295) );
  XNOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U339 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U340 ( .A(G106GAT), .B(KEYINPUT10), .Z(n299) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n307) );
  XNOR2_X1 U345 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n303), .B(G92GAT), .ZN(n342) );
  XOR2_X1 U347 ( .A(n342), .B(KEYINPUT67), .Z(n305) );
  XOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .Z(n443) );
  XNOR2_X1 U349 ( .A(n443), .B(G218GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U351 ( .A(n307), .B(n306), .Z(n311) );
  XNOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n308), .B(KEYINPUT7), .ZN(n385) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(G162GAT), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n309), .B(KEYINPUT78), .ZN(n425) );
  XNOR2_X1 U356 ( .A(n385), .B(n425), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n557) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n313) );
  XNOR2_X1 U359 ( .A(G57GAT), .B(G148GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n315) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n433) );
  XOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .Z(n439) );
  XOR2_X1 U365 ( .A(n433), .B(n439), .Z(n317) );
  XNOR2_X1 U366 ( .A(G29GAT), .B(G134GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n332) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT1), .Z(n321) );
  XNOR2_X1 U370 ( .A(G162GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U372 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n323) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G120GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U375 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n327) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U379 ( .A(G127GAT), .B(n328), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n518) );
  INV_X1 U382 ( .A(KEYINPUT33), .ZN(n333) );
  NAND2_X1 U383 ( .A1(KEYINPUT77), .A2(n333), .ZN(n336) );
  INV_X1 U384 ( .A(KEYINPUT77), .ZN(n334) );
  NAND2_X1 U385 ( .A1(n334), .A2(KEYINPUT33), .ZN(n335) );
  NAND2_X1 U386 ( .A1(n336), .A2(n335), .ZN(n338) );
  XNOR2_X1 U387 ( .A(KEYINPUT76), .B(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n340) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n339), .B(G64GAT), .ZN(n366) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G120GAT), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n341), .B(G71GAT), .ZN(n447) );
  XNOR2_X1 U393 ( .A(n447), .B(n342), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n291), .B(n343), .ZN(n346) );
  XOR2_X1 U395 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n345) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U397 ( .A(KEYINPUT73), .B(G204GAT), .Z(n348) );
  XNOR2_X1 U398 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U400 ( .A(G148GAT), .B(G106GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n436) );
  INV_X1 U402 ( .A(n436), .ZN(n351) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(n351), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(G211GAT), .Z(n355) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U407 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n357) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U410 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U411 ( .A(G78GAT), .B(G71GAT), .Z(n361) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(G8GAT), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(n362), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U417 ( .A(n365), .B(n428), .Z(n368) );
  XOR2_X1 U418 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XNOR2_X1 U419 ( .A(n440), .B(n366), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n582) );
  INV_X1 U421 ( .A(KEYINPUT36), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n557), .B(KEYINPUT105), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n586) );
  OR2_X1 U424 ( .A1(n582), .A2(n586), .ZN(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT45), .B(n371), .ZN(n372) );
  NOR2_X1 U426 ( .A1(n578), .A2(n372), .ZN(n390) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n374) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G1GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U430 ( .A(G197GAT), .B(KEYINPUT69), .Z(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n389) );
  XOR2_X1 U434 ( .A(G36GAT), .B(G8GAT), .Z(n415) );
  XOR2_X1 U435 ( .A(G113GAT), .B(G141GAT), .Z(n380) );
  XNOR2_X1 U436 ( .A(G43GAT), .B(G50GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(n415), .B(n381), .Z(n383) );
  NAND2_X1 U439 ( .A1(G229GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U441 ( .A(n384), .B(G15GAT), .Z(n387) );
  XNOR2_X1 U442 ( .A(n385), .B(G22GAT), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n572) );
  NAND2_X1 U445 ( .A1(n390), .A2(n572), .ZN(n399) );
  NAND2_X1 U446 ( .A1(n557), .A2(n582), .ZN(n394) );
  INV_X1 U447 ( .A(n572), .ZN(n533) );
  XOR2_X1 U448 ( .A(KEYINPUT41), .B(n578), .Z(n537) );
  NAND2_X1 U449 ( .A1(n533), .A2(n537), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U451 ( .A1(n394), .A2(n393), .ZN(n397) );
  INV_X1 U452 ( .A(KEYINPUT47), .ZN(n395) );
  NAND2_X1 U453 ( .A1(n399), .A2(n398), .ZN(n401) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n528) );
  INV_X1 U456 ( .A(n528), .ZN(n421) );
  XOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n403) );
  XNOR2_X1 U458 ( .A(G176GAT), .B(G183GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U460 ( .A(n404), .B(G190GAT), .Z(n406) );
  XNOR2_X1 U461 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n454) );
  XOR2_X1 U463 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n408) );
  XNOR2_X1 U464 ( .A(G204GAT), .B(KEYINPUT94), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n454), .B(n409), .ZN(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT21), .B(G211GAT), .Z(n411) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(G218GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n432) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(n432), .Z(n413) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U473 ( .A(n414), .B(G64GAT), .Z(n417) );
  XNOR2_X1 U474 ( .A(n415), .B(G92GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n461) );
  NAND2_X1 U477 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n422), .B(KEYINPUT54), .ZN(n423) );
  NOR2_X1 U479 ( .A1(n518), .A2(n423), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT64), .ZN(n571) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT24), .Z(n427) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n428), .B(KEYINPUT22), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n429), .B(KEYINPUT23), .ZN(n430) );
  XOR2_X1 U486 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n468) );
  NAND2_X1 U490 ( .A1(n571), .A2(n468), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U492 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U495 ( .A(n444), .B(n443), .Z(n452) );
  XOR2_X1 U496 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n446) );
  XNOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n447), .B(KEYINPUT85), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n448), .B(KEYINPUT83), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(n529) );
  NAND2_X1 U504 ( .A1(n455), .A2(n529), .ZN(n568) );
  NOR2_X1 U505 ( .A1(n557), .A2(n568), .ZN(n458) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n480) );
  NOR2_X1 U507 ( .A1(n572), .A2(n578), .ZN(n496) );
  NAND2_X1 U508 ( .A1(n529), .A2(n420), .ZN(n459) );
  NAND2_X1 U509 ( .A1(n468), .A2(n459), .ZN(n460) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n460), .ZN(n465) );
  XOR2_X1 U511 ( .A(n461), .B(KEYINPUT27), .Z(n471) );
  NOR2_X1 U512 ( .A1(n529), .A2(n468), .ZN(n462) );
  XNOR2_X1 U513 ( .A(n462), .B(KEYINPUT26), .ZN(n570) );
  NAND2_X1 U514 ( .A1(n471), .A2(n570), .ZN(n463) );
  XOR2_X1 U515 ( .A(KEYINPUT98), .B(n463), .Z(n464) );
  NOR2_X1 U516 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U517 ( .A1(n518), .A2(n466), .ZN(n467) );
  XNOR2_X1 U518 ( .A(n467), .B(KEYINPUT99), .ZN(n475) );
  XOR2_X1 U519 ( .A(n468), .B(KEYINPUT68), .Z(n469) );
  XNOR2_X1 U520 ( .A(KEYINPUT28), .B(n469), .ZN(n532) );
  XNOR2_X1 U521 ( .A(KEYINPUT88), .B(n529), .ZN(n470) );
  NOR2_X1 U522 ( .A1(n532), .A2(n470), .ZN(n473) );
  NAND2_X1 U523 ( .A1(n471), .A2(n518), .ZN(n472) );
  XNOR2_X1 U524 ( .A(n472), .B(KEYINPUT97), .ZN(n526) );
  NAND2_X1 U525 ( .A1(n473), .A2(n526), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n475), .A2(n474), .ZN(n492) );
  INV_X1 U527 ( .A(n582), .ZN(n541) );
  NAND2_X1 U528 ( .A1(n557), .A2(n541), .ZN(n476) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n476), .Z(n477) );
  AND2_X1 U530 ( .A1(n492), .A2(n477), .ZN(n505) );
  NAND2_X1 U531 ( .A1(n496), .A2(n505), .ZN(n478) );
  XOR2_X1 U532 ( .A(KEYINPUT100), .B(n478), .Z(n486) );
  NAND2_X1 U533 ( .A1(n518), .A2(n486), .ZN(n479) );
  XNOR2_X1 U534 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  XOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT101), .Z(n482) );
  NAND2_X1 U536 ( .A1(n486), .A2(n420), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n482), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n484) );
  NAND2_X1 U539 ( .A1(n486), .A2(n529), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT103), .Z(n488) );
  NAND2_X1 U543 ( .A1(n486), .A2(n532), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(n499) );
  XOR2_X1 U548 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n491), .ZN(n495) );
  NAND2_X1 U550 ( .A1(n582), .A2(n492), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n586), .A2(n493), .ZN(n494) );
  XOR2_X1 U552 ( .A(n495), .B(n494), .Z(n516) );
  NAND2_X1 U553 ( .A1(n516), .A2(n496), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n497), .Z(n503) );
  NAND2_X1 U555 ( .A1(n518), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n503), .A2(n420), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n503), .A2(n529), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n503), .A2(n532), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n507) );
  INV_X1 U565 ( .A(n537), .ZN(n562) );
  NOR2_X1 U566 ( .A1(n533), .A2(n562), .ZN(n515) );
  AND2_X1 U567 ( .A1(n515), .A2(n505), .ZN(n512) );
  NAND2_X1 U568 ( .A1(n512), .A2(n518), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n420), .A2(n512), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n529), .A2(n512), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U577 ( .A1(n512), .A2(n532), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(KEYINPUT111), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n420), .A2(n523), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n532), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n535) );
  INV_X1 U592 ( .A(n526), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n548) );
  NAND2_X1 U594 ( .A1(n548), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n530), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n545), .A2(n533), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U601 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  NAND2_X1 U604 ( .A1(n541), .A2(n545), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  INV_X1 U608 ( .A(n557), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n570), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n572), .A2(n556), .ZN(n549) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n549), .Z(n550) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U615 ( .A1(n556), .A2(n562), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n582), .A2(n556), .ZN(n555) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(n558), .Z(n559) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n572), .A2(n568), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n568), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n582), .A2(n568), .ZN(n569) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n585) );
  NOR2_X1 U637 ( .A1(n572), .A2(n585), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U644 ( .A(n585), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n583) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(n583), .Z(n584) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

