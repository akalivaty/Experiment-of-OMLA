//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n207), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n206), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n210), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n225), .B(new_n227), .C1(new_n218), .C2(new_n214), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n229));
  AND3_X1   g0029(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n230));
  AOI21_X1  g0030(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n229), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NOR3_X1   g0039(.A1(new_n222), .A2(new_n224), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(G361));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT68), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G250), .B(G257), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n263), .A3(G274), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n260), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n213), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G232), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n268), .B(new_n270), .C1(new_n207), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n262), .B1(new_n230), .B2(new_n231), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n266), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AND4_X1   g0086(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT73), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n259), .A2(G20), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n288), .A2(G77), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT15), .B(G87), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n284), .A2(G77), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n294), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n280), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n275), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n309), .B(new_n312), .C1(new_n313), .C2(new_n275), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G222), .A2(G1698), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n269), .A2(G223), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n267), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n273), .B(new_n318), .C1(G77), .C2(new_n267), .ZN(new_n319));
  INV_X1    g0119(.A(new_n265), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT70), .B(G226), .Z(new_n321));
  INV_X1    g0121(.A(G274), .ZN(new_n322));
  INV_X1    g0122(.A(new_n281), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n262), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n320), .A2(new_n321), .B1(new_n324), .B2(new_n261), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n276), .ZN(new_n327));
  OAI21_X1  g0127(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n328));
  INV_X1    g0128(.A(G150), .ZN(new_n329));
  INV_X1    g0129(.A(new_n299), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT8), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT71), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n202), .ZN(new_n334));
  NAND3_X1  g0134(.A1(KEYINPUT71), .A2(KEYINPUT8), .A3(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n233), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n295), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n287), .A2(G50), .A3(new_n292), .ZN(new_n340));
  INV_X1    g0140(.A(new_n284), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n201), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n319), .A2(new_n325), .A3(new_n278), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n327), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n339), .A2(KEYINPUT9), .A3(new_n340), .A4(new_n342), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n326), .A2(G200), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n319), .A2(new_n325), .A3(G190), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT10), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n347), .A4(new_n349), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n345), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n358));
  INV_X1    g0158(.A(G226), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n269), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n217), .A2(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n267), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n304), .B2(new_n206), .ZN(new_n364));
  NAND3_X1  g0164(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n273), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n320), .A2(G238), .B1(new_n324), .B2(new_n261), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n272), .B1(new_n362), .B2(new_n366), .ZN(new_n371));
  INV_X1    g0171(.A(G238), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n264), .B1(new_n265), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n358), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G169), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n371), .A2(new_n373), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT76), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT76), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(KEYINPUT13), .C1(new_n371), .C2(new_n373), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n358), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n380), .A2(G179), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(G169), .C1(new_n370), .C2(new_n375), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n377), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G68), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n305), .A2(G77), .B1(G20), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n201), .B2(new_n330), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT11), .B1(new_n390), .B2(new_n295), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n284), .A2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT77), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT12), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n394), .B(new_n395), .C1(KEYINPUT77), .C2(new_n392), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND4_X1   g0200(.A1(G68), .A2(new_n288), .A3(new_n291), .A4(new_n292), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n387), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n380), .A2(G190), .A3(new_n382), .A4(new_n383), .ZN(new_n405));
  OAI21_X1  g0205(.A(G200), .B1(new_n370), .B2(new_n375), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n315), .A2(new_n357), .A3(new_n404), .A4(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n202), .A2(new_n388), .ZN(new_n409));
  NOR2_X1   g0209(.A1(G58), .A2(G68), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n299), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G33), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n233), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(G20), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n419), .A2(new_n420), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT16), .B(new_n414), .C1(new_n422), .C2(new_n388), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT79), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n416), .A2(new_n417), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(KEYINPUT79), .A3(G33), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT80), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n416), .A2(new_n417), .A3(new_n424), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT80), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n421), .A4(new_n426), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n420), .B1(new_n267), .B2(G20), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n413), .B1(new_n433), .B2(G68), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n295), .B(new_n423), .C1(new_n434), .C2(KEYINPUT16), .ZN(new_n435));
  INV_X1    g0235(.A(new_n292), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n289), .A2(new_n336), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n341), .B2(new_n336), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n264), .B1(new_n265), .B2(new_n217), .ZN(new_n441));
  OR2_X1    g0241(.A1(G223), .A2(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n359), .A2(G1698), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n416), .A2(new_n442), .A3(new_n417), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G87), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n272), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n445), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n440), .B(new_n441), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n273), .A3(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(new_n441), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT82), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n276), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n278), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n439), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT18), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n435), .A2(new_n438), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n445), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT81), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(new_n272), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n440), .B1(new_n462), .B2(new_n441), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(KEYINPUT82), .A3(new_n453), .ZN(new_n464));
  AOI21_X1  g0264(.A(G200), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n462), .A2(G190), .A3(new_n441), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n459), .B(KEYINPUT17), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n435), .B(new_n438), .C1(new_n465), .C2(new_n466), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n439), .A2(new_n471), .A3(new_n455), .A4(new_n456), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n458), .A2(new_n467), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n408), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n263), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n263), .A2(G274), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n480), .A2(new_n218), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n418), .B2(new_n213), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n416), .A3(new_n417), .A4(G244), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n267), .A2(G250), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n269), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n273), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G169), .B1(new_n483), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n418), .A2(new_n225), .ZN(new_n494));
  OAI21_X1  g0294(.A(G1698), .B1(new_n494), .B2(new_n484), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n487), .A2(new_n488), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n485), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n482), .B1(new_n497), .B2(new_n273), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n493), .B1(new_n278), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT83), .B(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT6), .B1(new_n208), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n505), .A2(new_n233), .B1(new_n212), .B2(new_n330), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n433), .A2(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(KEYINPUT84), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n433), .A2(new_n509), .A3(G107), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n296), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n284), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n304), .A2(G1), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n287), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT85), .B1(new_n289), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n512), .B1(new_n518), .B2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n499), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n483), .A2(new_n492), .A3(new_n313), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n498), .B2(G200), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n433), .A2(new_n509), .A3(G107), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n509), .B1(new_n433), .B2(G107), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n524), .A2(new_n525), .A3(new_n506), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n519), .B(new_n523), .C1(new_n526), .C2(new_n296), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n500), .B2(new_n337), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(new_n233), .A3(G68), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n364), .A2(KEYINPUT19), .A3(new_n365), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n233), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G87), .A2(G107), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n500), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n296), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n516), .B2(new_n517), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n303), .A2(new_n284), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n372), .A2(new_n269), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n213), .A2(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n416), .A2(new_n543), .A3(new_n417), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n272), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n478), .A2(new_n322), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n225), .B1(new_n477), .B2(G1), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n263), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n546), .A2(new_n550), .A3(new_n313), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n543), .A2(new_n544), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n267), .B1(G33), .B2(G116), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(new_n272), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(G200), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n513), .B1(new_n287), .B2(new_n515), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n289), .A2(KEYINPUT85), .A3(new_n514), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n303), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n532), .A2(new_n233), .B1(new_n500), .B2(new_n534), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n529), .A2(new_n530), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n295), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n540), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n278), .B(new_n549), .C1(new_n553), .C2(new_n272), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n276), .B1(new_n546), .B2(new_n550), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n541), .A2(new_n555), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n521), .A2(new_n527), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n416), .A2(new_n417), .A3(new_n233), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n267), .A2(new_n571), .A3(new_n233), .A4(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n233), .A2(KEYINPUT23), .A3(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n207), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n207), .A3(G20), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(KEYINPUT86), .B1(new_n579), .B2(G20), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n573), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n573), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n295), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n284), .A2(G107), .ZN(new_n586));
  XOR2_X1   g0386(.A(new_n586), .B(KEYINPUT25), .Z(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n518), .B2(G107), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n416), .A2(new_n417), .A3(G250), .A4(new_n269), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n273), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n479), .A2(G264), .A3(new_n263), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT87), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n479), .A2(new_n481), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n476), .A2(new_n478), .B1(new_n323), .B2(new_n262), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT87), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(G264), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n593), .A2(new_n595), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G200), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n596), .B1(new_n592), .B2(new_n273), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n604), .A2(new_n313), .A3(new_n594), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n585), .B(new_n588), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n604), .A2(new_n594), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n607), .A2(new_n276), .B1(new_n601), .B2(new_n278), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n585), .A2(new_n588), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n514), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n288), .A2(new_n291), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n341), .A2(new_n612), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n233), .A2(G116), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n206), .A2(KEYINPUT83), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G97), .ZN(new_n620));
  AOI21_X1  g0420(.A(G33), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n488), .A2(new_n233), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n295), .B(new_n617), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n616), .B1(new_n232), .B2(new_n286), .ZN(new_n626));
  INV_X1    g0426(.A(new_n622), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n500), .B2(G33), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT20), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n614), .B(new_n615), .C1(new_n625), .C2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n476), .A2(new_n478), .ZN(new_n631));
  AOI22_X1  g0431(.A1(G270), .A2(new_n598), .B1(new_n631), .B2(new_n324), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n416), .A2(new_n417), .A3(G264), .A4(G1698), .ZN(new_n633));
  INV_X1    g0433(.A(G303), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n267), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n418), .A2(new_n218), .A3(G1698), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n273), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n276), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n637), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G200), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(new_n624), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n626), .A2(KEYINPUT20), .A3(new_n628), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n612), .B2(new_n341), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n632), .A2(new_n637), .A3(G190), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n643), .A2(new_n614), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n630), .A2(KEYINPUT21), .A3(new_n638), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n632), .A2(new_n637), .A3(G179), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n630), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n641), .A2(new_n648), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n475), .A2(new_n568), .A3(new_n611), .A4(new_n652), .ZN(G372));
  AND2_X1   g0453(.A1(new_n467), .A2(new_n470), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n404), .B1(new_n655), .B2(new_n311), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n458), .A2(new_n472), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n353), .A2(new_n356), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n345), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n607), .A2(new_n313), .B1(new_n601), .B2(new_n602), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n609), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n630), .A2(KEYINPUT21), .A3(new_n638), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT21), .B1(new_n630), .B2(new_n638), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n632), .A2(new_n637), .A3(G179), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n646), .B2(new_n614), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n668), .B2(new_n610), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n521), .A3(new_n527), .A4(new_n567), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n563), .ZN(new_n672));
  INV_X1    g0472(.A(new_n566), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n567), .B(new_n499), .C1(new_n511), .C2(new_n520), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n519), .B1(new_n526), .B2(new_n296), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .A3(new_n499), .A4(new_n567), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n674), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n474), .B1(new_n671), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n661), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n259), .A2(new_n233), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G213), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(KEYINPUT27), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G343), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n646), .B2(new_n614), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n652), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n641), .A2(new_n649), .A3(new_n651), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT88), .B1(new_n693), .B2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT88), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n696), .B(new_n697), .C1(new_n690), .C2(new_n692), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n610), .ZN(new_n702));
  INV_X1    g0502(.A(new_n688), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n609), .A2(new_n703), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n606), .A2(new_n610), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT89), .B1(new_n668), .B2(new_n703), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n691), .A2(new_n712), .A3(new_n688), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n714), .A2(new_n707), .B1(new_n702), .B2(new_n688), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n227), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n535), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(G1), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n235), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g0521(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n722));
  XNOR2_X1  g0522(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR4_X1   g0523(.A1(new_n568), .A2(new_n611), .A3(new_n652), .A4(new_n703), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n546), .A2(new_n550), .ZN(new_n725));
  AND4_X1   g0525(.A1(new_n725), .A2(new_n593), .A3(new_n595), .A4(new_n600), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n498), .A3(new_n650), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n498), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n725), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n601), .A3(new_n642), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n726), .A2(new_n498), .A3(new_n650), .A4(KEYINPUT30), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n703), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n697), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n703), .B1(new_n680), .B2(new_n670), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n742), .B1(new_n746), .B2(new_n744), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n741), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n723), .B1(new_n748), .B2(G1), .ZN(G364));
  AND2_X1   g0549(.A1(new_n233), .A2(G13), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n259), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n717), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n701), .B(new_n754), .C1(G330), .C2(new_n693), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n267), .A2(new_n226), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n226), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n254), .A2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n227), .A2(new_n267), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n477), .B2(new_n236), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n232), .B1(G20), .B2(new_n276), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n753), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n313), .A2(new_n602), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n233), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n538), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n233), .A2(new_n278), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n602), .A3(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n772), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n388), .B1(new_n780), .B2(new_n201), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n775), .B(new_n781), .C1(G77), .C2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n233), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n206), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n777), .A2(new_n313), .A3(G200), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n418), .B(new_n788), .C1(G58), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n773), .A2(new_n313), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT92), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G107), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n773), .A2(new_n782), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT32), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n785), .A2(new_n790), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  INV_X1    g0603(.A(G329), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n783), .A2(new_n803), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n789), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n780), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n805), .B(new_n808), .C1(G326), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n787), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G294), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n796), .A2(G283), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT94), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(KEYINPUT94), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n778), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n418), .B1(new_n774), .B2(new_n634), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n802), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n771), .B1(new_n821), .B2(new_n764), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n693), .B2(new_n769), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n755), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n826), .A2(new_n779), .B1(new_n806), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n267), .B(new_n828), .C1(G116), .C2(new_n784), .ZN(new_n829));
  INV_X1    g0629(.A(new_n788), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n796), .A2(G87), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n780), .A2(new_n634), .B1(new_n774), .B2(new_n207), .ZN(new_n832));
  INV_X1    g0632(.A(new_n798), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G311), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n778), .A2(G150), .B1(G159), .B2(new_n784), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT96), .B(G143), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n780), .C1(new_n806), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n267), .B1(new_n774), .B2(new_n201), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G132), .B2(new_n833), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n843), .B1(new_n202), .B2(new_n787), .C1(new_n388), .C2(new_n795), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n835), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n765), .A2(new_n767), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT95), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n845), .A2(new_n764), .B1(new_n212), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT99), .B1(new_n309), .B2(new_n688), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n307), .A2(new_n308), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n293), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n703), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT98), .B1(new_n280), .B2(new_n309), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT98), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n852), .A2(new_n857), .A3(new_n277), .A4(new_n279), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n314), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n310), .A2(new_n703), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n861), .B2(new_n767), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n753), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n742), .A2(new_n861), .ZN(new_n864));
  INV_X1    g0664(.A(new_n859), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n742), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n754), .B1(new_n867), .B2(new_n741), .ZN(new_n868));
  INV_X1    g0668(.A(new_n741), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n864), .B2(new_n866), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT100), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  INV_X1    g0673(.A(new_n505), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n234), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OAI211_X1 g0678(.A(new_n236), .B(G77), .C1(new_n202), .C2(new_n388), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n201), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n259), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n423), .A2(new_n295), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n418), .A2(new_n421), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n432), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G68), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n886), .B2(new_n414), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n438), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n455), .A2(new_n456), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n463), .A2(new_n464), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n466), .B1(new_n891), .B2(new_n602), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n889), .B(new_n890), .C1(new_n892), .C2(new_n439), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n687), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n468), .B2(new_n889), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n439), .A2(new_n687), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n457), .A2(new_n468), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n894), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n473), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(new_n900), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n889), .B1(new_n892), .B2(new_n439), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n893), .A3(new_n894), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n894), .B1(new_n658), .B2(new_n654), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n901), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n903), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n906), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n403), .A2(new_n703), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n404), .A2(new_n407), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n403), .B(new_n703), .C1(new_n655), .C2(new_n387), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(new_n859), .B2(new_n860), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(KEYINPUT104), .C1(new_n724), .C2(new_n739), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n521), .A2(new_n527), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n611), .A2(new_n652), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n567), .A4(new_n688), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n737), .A3(new_n738), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT104), .B1(new_n926), .B2(new_n920), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT40), .B1(new_n916), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n899), .B1(new_n658), .B2(new_n654), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n457), .A2(new_n468), .A3(new_n899), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n932), .A2(new_n900), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n907), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n904), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n926), .A2(new_n920), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT40), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n929), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n475), .A2(new_n740), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n697), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n658), .A2(new_n687), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n703), .B1(new_n856), .B2(new_n858), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n742), .B2(new_n865), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n918), .A2(new_n919), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT101), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT101), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n703), .B(new_n859), .C1(new_n680), .C2(new_n670), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n946), .C1(new_n950), .C2(new_n944), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n915), .A2(new_n914), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n897), .A2(new_n900), .B1(new_n473), .B2(new_n902), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT103), .B1(new_n953), .B2(KEYINPUT38), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n948), .B(new_n951), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT39), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n904), .A2(new_n934), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n916), .B2(KEYINPUT39), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n387), .A2(new_n403), .A3(new_n688), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n943), .B(new_n955), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n745), .A2(new_n474), .A3(new_n747), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n661), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n942), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n259), .B2(new_n750), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n942), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n882), .B1(new_n965), .B2(new_n966), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n250), .A2(new_n760), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n770), .B1(new_n227), .B2(new_n303), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n754), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n779), .A2(new_n827), .B1(new_n780), .B2(new_n803), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n806), .A2(new_n634), .B1(new_n783), .B2(new_n826), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n267), .B1(new_n833), .B2(G317), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n207), .B2(new_n787), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n774), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT109), .B1(new_n976), .B2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n978), .C1(new_n500), .C2(new_n795), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n787), .A2(new_n388), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n418), .B(new_n980), .C1(G58), .C2(new_n976), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n796), .A2(G77), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n780), .A2(new_n838), .B1(new_n798), .B2(new_n837), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G150), .B2(new_n789), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n778), .A2(G159), .B1(G50), .B2(new_n784), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT110), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n979), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  OR2_X1    g0789(.A1(new_n541), .A2(new_n688), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT105), .Z(new_n991));
  MUX2_X1   g0791(.A(new_n674), .B(new_n567), .S(new_n991), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n970), .B1(new_n989), .B2(new_n765), .C1(new_n992), .C2(new_n769), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n751), .B(KEYINPUT108), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n694), .A2(new_n698), .A3(KEYINPUT106), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT106), .B1(new_n694), .B2(new_n698), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n714), .A2(new_n707), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n708), .A2(new_n713), .A3(new_n711), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n998), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n700), .A2(KEYINPUT106), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(KEYINPUT107), .A3(new_n748), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n678), .A2(new_n703), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n923), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n678), .A2(new_n499), .A3(new_n703), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n715), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT45), .Z(new_n1010));
  NOR2_X1   g0810(.A1(new_n715), .A2(new_n1008), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT44), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n709), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n710), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1004), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT107), .B1(new_n1003), .B2(new_n748), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n748), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n717), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n995), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1008), .A2(new_n707), .A3(new_n714), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n923), .A2(new_n702), .A3(new_n1005), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n703), .B1(new_n1024), .B2(new_n521), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1022), .B2(KEYINPUT42), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1023), .A2(new_n1026), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n1027), .A2(KEYINPUT43), .A3(new_n992), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n709), .A2(new_n1008), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n993), .B1(new_n1021), .B2(new_n1035), .ZN(G387));
  OR2_X1    g0836(.A1(new_n1003), .A2(new_n748), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1003), .A2(new_n748), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n717), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n708), .A2(new_n768), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n719), .A2(new_n756), .B1(G107), .B2(new_n226), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n298), .A2(new_n300), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n201), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT50), .Z(new_n1044));
  OAI211_X1 g0844(.A(new_n719), .B(new_n477), .C1(new_n388), .C2(new_n212), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT111), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n761), .B1(new_n246), .B2(G45), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n753), .B1(new_n1049), .B2(new_n770), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n774), .A2(new_n212), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n780), .A2(new_n799), .B1(new_n798), .B2(new_n329), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G50), .C2(new_n789), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n787), .A2(new_n302), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n418), .B(new_n1054), .C1(G68), .C2(new_n784), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n796), .A2(G97), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n778), .A2(new_n334), .A3(new_n335), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n780), .A2(new_n807), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n779), .A2(new_n803), .B1(new_n783), .B2(new_n634), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G317), .C2(new_n789), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(KEYINPUT48), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(KEYINPUT48), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n787), .A2(new_n826), .B1(new_n774), .B2(new_n827), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n796), .A2(G116), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n267), .B1(new_n833), .B2(G326), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1058), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1050), .B1(new_n1071), .B2(new_n764), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1003), .A2(new_n995), .B1(new_n1040), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1039), .A2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1017), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(new_n1004), .A3(new_n1015), .A4(new_n1014), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(new_n1014), .Z(new_n1078));
  INV_X1    g0878(.A(new_n1038), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n717), .B(new_n1076), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1006), .A2(new_n768), .A3(new_n1007), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n267), .B1(new_n774), .B2(new_n388), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n779), .A2(new_n201), .B1(new_n798), .B2(new_n838), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G77), .C2(new_n811), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n789), .A2(G159), .B1(new_n809), .B2(G150), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1042), .A2(new_n784), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n831), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n789), .A2(G311), .B1(new_n809), .B2(G317), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n779), .A2(new_n634), .B1(new_n783), .B2(new_n827), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G283), .B2(new_n976), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n418), .B1(new_n798), .B2(new_n807), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n811), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n797), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n765), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n257), .A2(new_n760), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n500), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n770), .B1(new_n227), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n754), .B(new_n1097), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT114), .Z(new_n1102));
  AOI22_X1  g0902(.A1(new_n1078), .A2(new_n995), .B1(new_n1081), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1080), .A2(new_n1103), .ZN(G390));
  OAI21_X1  g0904(.A(KEYINPUT39), .B1(new_n952), .B2(new_n954), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n944), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n866), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n946), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n959), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n957), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n959), .A3(new_n935), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n741), .A2(new_n861), .A3(new_n946), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1114), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n741), .A2(new_n474), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n961), .A2(new_n661), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n926), .A2(new_n861), .A3(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n947), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1107), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1114), .A2(new_n945), .A3(new_n1121), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1116), .A2(new_n1117), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT115), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1125), .B(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1111), .A2(new_n1114), .A3(new_n1112), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n717), .B(new_n1126), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n995), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n958), .A2(new_n766), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G107), .A2(new_n778), .B1(new_n789), .B2(G116), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n500), .B2(new_n783), .C1(new_n795), .C2(new_n388), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n809), .A2(G283), .B1(new_n833), .B2(G294), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n775), .A2(new_n267), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n212), .C2(new_n787), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n811), .A2(G159), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n329), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n418), .B1(new_n833), .B2(G125), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT53), .B1(new_n774), .B2(new_n329), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n778), .A2(G137), .B1(new_n809), .B2(G128), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n789), .A2(G132), .B1(new_n784), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(new_n1149), .C1(new_n795), .C2(new_n201), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1137), .A2(new_n1140), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n764), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n754), .B1(new_n848), .B2(new_n336), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1135), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1133), .A2(new_n1134), .A3(new_n1154), .ZN(G378));
  NOR2_X1   g0955(.A1(new_n357), .A2(KEYINPUT117), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n343), .A2(new_n687), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT118), .Z(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT117), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n345), .C1(new_n353), .C2(new_n356), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1157), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1159), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1169), .A2(KEYINPUT119), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT119), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n766), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n753), .B1(new_n846), .B2(G50), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT116), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n780), .A2(new_n1177), .B1(new_n783), .B2(new_n837), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n789), .A2(G128), .B1(new_n976), .B2(new_n1148), .ZN(new_n1179));
  INV_X1    g0979(.A(G132), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n779), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(G150), .C2(new_n811), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n796), .A2(G159), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n833), .C2(G124), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n796), .A2(G58), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n778), .A2(G97), .B1(G283), .B2(new_n833), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n302), .C2(new_n783), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n267), .A2(G41), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(new_n1051), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n806), .A2(new_n207), .B1(new_n780), .B2(new_n612), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1191), .A2(new_n980), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1192), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1195), .A2(KEYINPUT58), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1188), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1176), .B1(new_n1199), .B2(new_n764), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1174), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1169), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1170), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n904), .A2(new_n934), .ZN(new_n1207));
  OAI21_X1  g1007(.A(G330), .B1(new_n1207), .B2(new_n937), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n929), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n928), .B1(new_n952), .B2(new_n954), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT40), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n697), .B1(new_n938), .B2(new_n935), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(KEYINPUT120), .A3(new_n960), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n959), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n955), .A2(new_n943), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT120), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1209), .A3(new_n1215), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1202), .B1(new_n1222), .B2(new_n995), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1119), .B1(new_n1132), .B2(new_n1125), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n929), .A2(new_n1208), .A3(new_n1173), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1205), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n960), .A2(new_n1209), .A3(new_n1215), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(KEYINPUT57), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n717), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT121), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1119), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1126), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1222), .A2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1232), .A2(new_n1233), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(KEYINPUT121), .B(new_n717), .C1(new_n1225), .C2(new_n1231), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1224), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT122), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(G375));
  AOI21_X1  g1042(.A(new_n754), .B1(new_n848), .B2(new_n388), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n779), .A2(new_n1147), .B1(new_n783), .B2(new_n329), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n418), .B(new_n1244), .C1(G137), .C2(new_n789), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n811), .A2(G50), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n780), .A2(new_n1180), .B1(new_n774), .B2(new_n799), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G128), .B2(new_n833), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1189), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n774), .A2(new_n206), .B1(new_n798), .B2(new_n634), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n779), .A2(new_n612), .B1(new_n783), .B2(new_n207), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G283), .B2(new_n789), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n267), .B(new_n1054), .C1(G294), .C2(new_n809), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n982), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1251), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n764), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1243), .B1(new_n946), .B2(new_n767), .C1(new_n1257), .C2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(new_n994), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1123), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1020), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1129), .B2(new_n1265), .ZN(G381));
  INV_X1    g1066(.A(G387), .ZN(new_n1267));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1039), .A2(new_n824), .A3(new_n1073), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1241), .A2(new_n1267), .A3(new_n1268), .A4(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n1241), .A2(new_n1268), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1269), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(G387), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1019), .B1(new_n1076), .B2(new_n748), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1034), .B1(new_n1280), .B2(new_n995), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1276), .B1(new_n1281), .B2(new_n993), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1274), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1277), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1281), .B2(new_n993), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1284), .B(G390), .C1(new_n1285), .C2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1264), .B1(new_n1125), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1261), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n717), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1291), .A3(new_n1294), .A4(new_n717), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1296), .B2(new_n1263), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n872), .B(new_n1262), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G343), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(G213), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(G2897), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G2897), .B(new_n1302), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1222), .A2(new_n1236), .A3(new_n1020), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1202), .B1(new_n1308), .B2(new_n995), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G378), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1240), .B2(G378), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1306), .B1(new_n1311), .B2(new_n1302), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1216), .B(new_n1220), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1234), .B1(new_n1313), .B2(new_n1225), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1229), .A2(KEYINPUT57), .A3(new_n1230), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n718), .B1(new_n1315), .B2(new_n1236), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1316), .B2(KEYINPUT121), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1239), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1223), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1309), .A2(new_n1307), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1268), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1301), .A4(new_n1299), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1312), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1302), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1323), .B1(new_n1327), .B2(new_n1299), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1288), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1299), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1333), .B1(new_n1287), .B2(new_n1325), .ZN(new_n1334));
  AOI211_X1 g1134(.A(KEYINPUT127), .B(KEYINPUT61), .C1(new_n1283), .C2(new_n1286), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1327), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1332), .A2(new_n1336), .A3(new_n1312), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1329), .A2(new_n1338), .ZN(G405));
  OR2_X1    g1139(.A1(new_n1240), .A2(new_n1268), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1272), .A2(new_n1340), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1287), .B(new_n1299), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1272), .A3(new_n1340), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(G402));
endmodule


