//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n447, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(G137), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XOR2_X1   g054(.A(KEYINPUT3), .B(G2104), .Z(new_n480));
  OR3_X1    g055(.A1(new_n480), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n480), .B2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT68), .Z(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n473), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n480), .A2(new_n476), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n486), .A2(new_n488), .B1(new_n489), .B2(G124), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n484), .A2(new_n490), .ZN(G162));
  AND3_X1   g066(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n492));
  AND2_X1   g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n476), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n467), .A2(G126), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n467), .B(KEYINPUT66), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G138), .A3(new_n476), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n505), .B2(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n515), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT69), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n505), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  OAI211_X1 g096(.A(G543), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(new_n521), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n518), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n505), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n537), .B1(new_n513), .B2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n515), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(new_n539), .B1(new_n513), .B2(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n540), .A2(KEYINPUT72), .A3(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n534), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n533), .A2(new_n542), .ZN(G168));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n536), .B2(new_n541), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n540), .A2(new_n505), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n515), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n536), .B2(new_n541), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n546), .A2(new_n553), .B1(new_n554), .B2(new_n515), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT73), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT73), .B1(new_n552), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(G65), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n505), .A2(new_n566), .B1(G78), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n515), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(new_n570), .B1(G91), .B2(new_n520), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n522), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n540), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(KEYINPUT74), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n571), .A2(new_n578), .A3(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  NAND2_X1  g157(.A1(new_n520), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n523), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n520), .A2(G86), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n505), .A2(KEYINPUT77), .A3(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(KEYINPUT77), .B1(new_n505), .B2(G61), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n536), .A2(new_n541), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n597), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n546), .A2(new_n599), .B1(new_n600), .B2(new_n515), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n598), .A2(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n520), .A2(G92), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n522), .A2(new_n535), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT72), .B1(new_n540), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT79), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n536), .A2(new_n541), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n607), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n505), .A2(G66), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT80), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n515), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n536), .A2(new_n611), .A3(new_n541), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n611), .B1(new_n536), .B2(new_n541), .ZN(new_n620));
  OAI21_X1  g195(.A(G54), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  INV_X1    g197(.A(new_n617), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n606), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n604), .B1(new_n625), .B2(new_n603), .ZN(G284));
  AOI21_X1  g201(.A(new_n604), .B1(new_n625), .B2(new_n603), .ZN(G321));
  MUX2_X1   g202(.A(G286), .B(G299), .S(new_n603), .Z(G280));
  XNOR2_X1  g203(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n625), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n559), .A2(new_n603), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n630), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n603), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n483), .A2(G135), .ZN(new_n637));
  MUX2_X1   g212(.A(G99), .B(G111), .S(G2105), .Z(new_n638));
  AOI22_X1  g213(.A1(new_n489), .A2(G123), .B1(G2104), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT85), .B(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n499), .A2(new_n474), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT13), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2427), .ZN(new_n652));
  INV_X1    g227(.A(G2430), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(KEYINPUT17), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n666), .A3(new_n668), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n668), .B1(new_n666), .B2(new_n667), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n674), .A2(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(KEYINPUT87), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n666), .B2(new_n672), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n671), .B(new_n673), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G2096), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(G227));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n687), .A3(new_n685), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n692), .C1(new_n687), .C2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT32), .B(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1971), .Z(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT33), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT34), .B1(new_n705), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n705), .A2(new_n715), .A3(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G24), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n598), .A2(new_n601), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT89), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n719), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1986), .ZN(new_n723));
  NOR2_X1   g298(.A1(G25), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n483), .A2(G131), .ZN(new_n725));
  MUX2_X1   g300(.A(G95), .B(G107), .S(G2105), .Z(new_n726));
  AOI22_X1  g301(.A1(new_n489), .A2(G119), .B1(G2104), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  NOR3_X1   g307(.A1(new_n718), .A2(new_n723), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n717), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT36), .ZN(new_n735));
  NOR2_X1   g310(.A1(G168), .A2(new_n709), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n709), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G35), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G162), .B2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n739), .B1(new_n742), .B2(G2090), .ZN(new_n743));
  NOR2_X1   g318(.A1(G27), .A2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G164), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(new_n443), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n483), .A2(G141), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n474), .A2(G105), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G129), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G32), .B(new_n756), .S(G29), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n640), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT30), .A2(G28), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT30), .A2(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT31), .B(G11), .Z(new_n765));
  NOR3_X1   g340(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n746), .A2(new_n759), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n760), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n481), .A2(G140), .A3(new_n482), .ZN(new_n770));
  MUX2_X1   g345(.A(G104), .B(G116), .S(G2105), .Z(new_n771));
  AOI22_X1  g346(.A1(new_n489), .A2(G128), .B1(G2104), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n769), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G160), .B2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(G2084), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n743), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n709), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n559), .B2(new_n709), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1341), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n709), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n709), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n709), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G1961), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1961), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n737), .B2(new_n738), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n792), .B(new_n794), .C1(new_n742), .C2(G2090), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n782), .A2(new_n785), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n625), .B2(G16), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1348), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(G1348), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n760), .A2(G33), .ZN(new_n802));
  NAND2_X1  g377(.A1(G115), .A2(G2104), .ZN(new_n803));
  INV_X1    g378(.A(G127), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n469), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n805), .A2(KEYINPUT92), .A3(G2105), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT92), .B1(new_n805), .B2(G2105), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n474), .A2(G103), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n481), .A2(new_n482), .ZN(new_n811));
  INV_X1    g386(.A(G139), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n806), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n802), .B1(new_n815), .B2(G29), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n442), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n780), .A2(G2084), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n757), .B2(new_n758), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n816), .B2(new_n442), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(KEYINPUT96), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n801), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT96), .B1(new_n818), .B2(new_n821), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n735), .A2(new_n825), .ZN(G150));
  XNOR2_X1  g401(.A(G150), .B(KEYINPUT97), .ZN(G311));
  INV_X1    g402(.A(new_n606), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n617), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n630), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n597), .A2(G55), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n519), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n520), .A2(G93), .B1(new_n837), .B2(G651), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n556), .A2(new_n557), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n834), .B(new_n838), .C1(new_n552), .C2(new_n555), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n833), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n839), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT98), .ZN(G145));
  NOR2_X1   g425(.A1(new_n756), .A2(new_n773), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n770), .A2(new_n772), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n747), .B2(new_n755), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n498), .A2(new_n502), .A3(KEYINPUT99), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT99), .B1(new_n498), .B2(new_n502), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n851), .A2(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n756), .A2(new_n773), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n747), .A3(new_n755), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n503), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n854), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT100), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n814), .B1(new_n863), .B2(KEYINPUT93), .ZN(new_n864));
  INV_X1    g439(.A(new_n814), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n857), .A3(new_n862), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  MUX2_X1   g447(.A(G106), .B(G118), .S(G2105), .Z(new_n873));
  AOI22_X1  g448(.A1(new_n489), .A2(G130), .B1(G2104), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G142), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n811), .B2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n645), .B(new_n876), .Z(new_n877));
  NAND3_X1  g452(.A1(new_n725), .A2(KEYINPUT101), .A3(new_n727), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT101), .B1(new_n725), .B2(new_n727), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n728), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT102), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n877), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n645), .B(new_n876), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(KEYINPUT102), .A3(new_n878), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n872), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n872), .A3(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n871), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n886), .A2(new_n872), .A3(new_n890), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n864), .B(new_n870), .C1(new_n895), .C2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G162), .B(new_n478), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n640), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n640), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n886), .A2(new_n890), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT104), .B1(new_n864), .B2(new_n870), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT106), .B1(new_n900), .B2(new_n901), .ZN(new_n909));
  INV_X1    g484(.A(new_n901), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n899), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n895), .A2(new_n891), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n871), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(new_n862), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n858), .A2(new_n859), .B1(new_n861), .B2(new_n854), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n865), .B1(new_n920), .B2(new_n866), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n869), .A2(new_n857), .A3(new_n862), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n904), .B1(new_n925), .B2(new_n905), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n903), .B1(new_n916), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g503(.A1(new_n839), .A2(G868), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n633), .B(new_n842), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  INV_X1    g506(.A(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n618), .A2(new_n624), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n828), .ZN(new_n934));
  AOI211_X1 g509(.A(G299), .B(new_n606), .C1(new_n618), .C2(new_n624), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n831), .A2(G299), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n625), .A2(new_n932), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  XOR2_X1   g518(.A(G303), .B(KEYINPUT107), .Z(new_n944));
  AND2_X1   g519(.A1(new_n944), .A2(new_n702), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n702), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n720), .B(new_n711), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n943), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n929), .B1(new_n951), .B2(G868), .ZN(G295));
  AOI21_X1  g527(.A(new_n929), .B1(new_n951), .B2(G868), .ZN(G331));
  INV_X1    g528(.A(new_n542), .ZN(new_n954));
  INV_X1    g529(.A(new_n532), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n529), .B2(new_n505), .ZN(new_n956));
  NAND3_X1  g531(.A1(G171), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n533), .A2(new_n542), .B1(new_n545), .B2(new_n549), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n959), .A2(new_n840), .A3(new_n841), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n841), .B2(new_n840), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n936), .A2(new_n939), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n937), .A3(new_n938), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(KEYINPUT108), .A3(new_n965), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n950), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n950), .A2(new_n963), .A3(new_n965), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n950), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n963), .A2(KEYINPUT108), .A3(new_n965), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT108), .B1(new_n963), .B2(new_n965), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n971), .A2(new_n972), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n963), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n936), .A2(new_n939), .A3(new_n962), .A4(KEYINPUT110), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n965), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n964), .A2(KEYINPUT111), .A3(new_n937), .A4(new_n938), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n986), .A2(new_n987), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n973), .B1(new_n991), .B2(new_n977), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n986), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n977), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND4_X1   g572(.A1(new_n984), .A2(new_n997), .A3(new_n993), .A4(new_n981), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n976), .B(new_n983), .C1(new_n994), .C2(new_n998), .ZN(new_n999));
  MUX2_X1   g574(.A(new_n992), .B(new_n982), .S(new_n993), .Z(new_n1000));
  MUX2_X1   g575(.A(new_n999), .B(new_n1000), .S(KEYINPUT44), .Z(G397));
  XOR2_X1   g576(.A(KEYINPUT113), .B(G40), .Z(new_n1002));
  OR2_X1    g577(.A1(new_n478), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n503), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT48), .Z(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n756), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n852), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n773), .A2(G2067), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n728), .B(new_n731), .Z(new_n1019));
  OAI21_X1  g594(.A(new_n1008), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1011), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1009), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1008), .A2(KEYINPUT125), .A3(KEYINPUT46), .A4(new_n1012), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1017), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1008), .B1(new_n756), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n729), .A2(new_n731), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1030), .B(KEYINPUT124), .Z(new_n1031));
  OAI21_X1  g606(.A(new_n1015), .B1(new_n1031), .B2(new_n1018), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1008), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1021), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT126), .ZN(new_n1035));
  OR2_X1    g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n595), .A2(new_n587), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G1981), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT115), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n711), .B2(G1976), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(G1976), .B2(new_n711), .ZN(new_n1048));
  MUX2_X1   g623(.A(new_n1046), .B(new_n1047), .S(new_n1048), .Z(new_n1049));
  AND2_X1   g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n478), .A2(new_n1002), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT45), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1007), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1054), .A2(G1971), .B1(new_n1058), .B2(G2090), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G303), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT55), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1007), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n738), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n1051), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1068), .A2(G8), .A3(G168), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1063), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1050), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1036), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1045), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1045), .A2(new_n1049), .A3(new_n1069), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1060), .B(KEYINPUT116), .Z(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1062), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g655(.A(new_n1074), .B1(new_n1077), .B2(new_n1043), .C1(new_n1080), .C2(new_n1070), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(G8), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT121), .Z(new_n1083));
  AOI211_X1 g658(.A(KEYINPUT51), .B(new_n1083), .C1(new_n1068), .C2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1007), .A2(new_n443), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1058), .A2(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  XOR2_X1   g664(.A(G171), .B(KEYINPUT54), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT122), .B(G2078), .ZN(new_n1092));
  NAND2_X1  g667(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n478), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1007), .A3(new_n1053), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT123), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1088), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1065), .A2(new_n1101), .A3(new_n1067), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(G8), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1083), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1083), .A3(new_n1102), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(KEYINPUT51), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1084), .B(new_n1099), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1054), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1054), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1058), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1111), .B(new_n1113), .C1(G1956), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n571), .A2(new_n576), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT61), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(new_n1125), .B1(new_n1064), .B2(G1996), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n559), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1058), .A2(new_n1129), .B1(new_n1124), .B2(new_n1014), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(new_n831), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n831), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(new_n1134), .A3(new_n625), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1128), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1122), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1120), .B(KEYINPUT119), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1115), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1122), .A2(KEYINPUT61), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1108), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1089), .A2(G171), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1084), .B1(new_n1107), .B2(new_n1105), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT62), .B(new_n1084), .C1(new_n1107), .C2(new_n1105), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1050), .A2(new_n1072), .A3(new_n1063), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1081), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G290), .B(G1986), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1008), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT114), .Z(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1020), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1035), .B1(new_n1153), .B2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g733(.A1(G229), .A2(new_n464), .A3(G401), .A4(G227), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n927), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g735(.A(KEYINPUT109), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n1162));
  AOI211_X1 g736(.A(new_n975), .B(new_n993), .C1(new_n980), .C2(new_n981), .ZN(new_n1163));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n997), .A2(new_n993), .A3(new_n981), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1165), .A2(KEYINPUT112), .ZN(new_n1166));
  NAND3_X1  g740(.A1(new_n992), .A2(new_n984), .A3(new_n993), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g742(.A(KEYINPUT127), .B(new_n1161), .C1(new_n1164), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  INV_X1    g744(.A(new_n1161), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n999), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1169), .A2(new_n1172), .ZN(G308));
  NAND2_X1  g747(.A1(new_n999), .A2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n999), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1176), .ZN(G225));
endmodule


