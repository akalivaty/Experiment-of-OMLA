//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n210), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(G244), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n217), .A2(G77), .B1(KEYINPUT65), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n218), .C2(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n216), .B(new_n227), .C1(KEYINPUT0), .C2(new_n210), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT13), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  AND3_X1   g0049(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(new_n246), .B2(new_n248), .ZN(new_n251));
  OAI211_X1 g0051(.A(G232), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  OAI211_X1 g0053(.A(G226), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G41), .A2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n263), .A3(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT67), .A2(G1), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT67), .A2(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n267), .B2(new_n261), .ZN(new_n268));
  INV_X1    g0068(.A(G238), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n244), .B1(new_n260), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI211_X1 g0073(.A(KEYINPUT13), .B(new_n270), .C1(new_n256), .C2(new_n259), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G190), .ZN(new_n276));
  OAI21_X1  g0076(.A(G200), .B1(new_n272), .B2(new_n274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n212), .A2(G33), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n279), .B1(new_n212), .B2(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n211), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(KEYINPUT11), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(KEYINPUT11), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n283), .A2(new_n211), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n267), .B2(new_n212), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(G13), .B(G20), .C1(new_n265), .C2(new_n266), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G68), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n276), .A2(new_n277), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n272), .A2(new_n274), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT14), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(G169), .C1(new_n272), .C2(new_n274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(G179), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n295), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n264), .B1(new_n268), .B2(new_n224), .ZN(new_n307));
  OAI211_X1 g0107(.A(G222), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n308));
  OAI211_X1 g0108(.A(G223), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n247), .A2(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT68), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G77), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n308), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n307), .B1(new_n315), .B2(new_n259), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G190), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT8), .A2(G58), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT8), .A2(G58), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n281), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n322), .B1(G150), .B2(new_n278), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n203), .A2(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n289), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT67), .B(G1), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n326), .A2(G13), .A3(G20), .A4(new_n202), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n290), .B2(new_n202), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n318), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n278), .A2(G150), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n319), .A2(new_n320), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n324), .B(new_n330), .C1(new_n331), .C2(new_n281), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n284), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n284), .B1(new_n326), .B2(G20), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G50), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(KEYINPUT9), .A3(new_n327), .A4(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n317), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n316), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT10), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n316), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n317), .A4(new_n337), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(G238), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n347));
  INV_X1    g0147(.A(G107), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n312), .A2(new_n313), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n349), .A2(G232), .A3(new_n253), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n259), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n217), .B(new_n258), .C1(new_n267), .C2(new_n261), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n353), .A2(KEYINPUT69), .A3(new_n264), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT69), .B1(new_n353), .B2(new_n264), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n356), .A3(G190), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n290), .A2(new_n280), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n321), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n359));
  OR2_X1    g0159(.A1(KEYINPUT15), .A2(G87), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT15), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n322), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n289), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n292), .ZN(new_n364));
  AOI211_X1 g0164(.A(new_n358), .B(new_n363), .C1(new_n280), .C2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n352), .A2(new_n356), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n367), .B2(new_n298), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n352), .A2(new_n356), .A3(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n366), .A2(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n342), .A2(G179), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n333), .A2(new_n327), .A3(new_n335), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n316), .B2(G169), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AND4_X1   g0177(.A1(new_n306), .A2(new_n346), .A3(new_n372), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n341), .B2(new_n345), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n306), .B1(new_n379), .B2(new_n372), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n305), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(G232), .B(new_n258), .C1(new_n267), .C2(new_n261), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G223), .A2(G1698), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n224), .B2(G1698), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT3), .B(G33), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(G33), .B2(G87), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n382), .B(new_n264), .C1(new_n386), .C2(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G169), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n370), .B2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n385), .A2(new_n390), .A3(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n246), .A2(new_n248), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(new_n212), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G58), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n288), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n201), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n278), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n284), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n312), .A2(new_n212), .A3(new_n313), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n391), .B1(new_n404), .B2(new_n390), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(new_n288), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n292), .A2(new_n331), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n334), .B2(new_n331), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT18), .B(new_n389), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n403), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n390), .B1(new_n385), .B2(G20), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n399), .B1(new_n418), .B2(G68), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n289), .B1(new_n419), .B2(KEYINPUT16), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT72), .A3(KEYINPUT18), .A4(new_n389), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  INV_X1    g0224(.A(new_n389), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n414), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n415), .A2(new_n420), .ZN(new_n428));
  INV_X1    g0228(.A(new_n411), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n387), .A2(G200), .ZN(new_n430));
  INV_X1    g0230(.A(new_n264), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n224), .A2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G223), .B2(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n433), .A2(new_n392), .B1(new_n245), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n431), .B1(new_n435), .B2(new_n259), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G190), .A3(new_n382), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n429), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n427), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n381), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT4), .ZN(new_n446));
  INV_X1    g0246(.A(G244), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n253), .B(new_n448), .C1(new_n250), .C2(new_n251), .ZN(new_n449));
  OAI211_X1 g0249(.A(G250), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n246), .A2(new_n248), .A3(G244), .A4(new_n253), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n446), .B1(G33), .B2(G283), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n259), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT74), .B1(new_n455), .B2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT74), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(G41), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n258), .A2(G274), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT75), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  INV_X1    g0264(.A(new_n266), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT67), .A2(G1), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n326), .A2(G45), .A3(G274), .A4(new_n258), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT75), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n259), .B1(new_n461), .B2(new_n467), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n468), .A2(new_n471), .B1(new_n472), .B2(G257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n454), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n364), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G33), .B1(new_n265), .B2(new_n266), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n292), .A2(new_n289), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(new_n476), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n348), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n238), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(KEYINPUT6), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n405), .B2(new_n348), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n480), .B1(new_n485), .B2(new_n284), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n454), .A2(G190), .A3(new_n473), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n454), .A2(new_n370), .A3(new_n473), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(G169), .B1(new_n454), .B2(new_n473), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n490), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT76), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n486), .A2(new_n491), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n489), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT78), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n250), .A2(new_n251), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G257), .A2(G1698), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n253), .A2(G264), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n392), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n259), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n471), .A2(new_n468), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n472), .A2(G270), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n292), .A2(new_n478), .A3(G116), .A4(new_n289), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n326), .A2(G13), .A3(G20), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n283), .A2(new_n211), .B1(G20), .B2(new_n512), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(G33), .B2(G283), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G33), .B2(new_n476), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n298), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n501), .B1(new_n510), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT78), .B1(new_n510), .B2(new_n523), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n500), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n510), .A2(new_n523), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT78), .B(KEYINPUT21), .C1(new_n528), .C2(new_n501), .ZN(new_n529));
  AND4_X1   g0329(.A1(G179), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n514), .A2(new_n522), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n510), .B2(G200), .ZN(new_n533));
  INV_X1    g0333(.A(G190), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n510), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n527), .A2(new_n529), .A3(new_n532), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n269), .A2(new_n253), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n447), .A2(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n246), .A2(new_n537), .A3(new_n248), .A4(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n245), .A2(new_n512), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n259), .ZN(new_n543));
  OAI21_X1  g0343(.A(G45), .B1(new_n265), .B2(new_n266), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(G250), .A3(new_n258), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n543), .A2(G190), .A3(new_n469), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n469), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n258), .B1(new_n539), .B2(new_n541), .ZN(new_n548));
  OAI21_X1  g0348(.A(G200), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n479), .A2(new_n434), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n212), .B1(new_n255), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n434), .A2(new_n476), .A3(new_n348), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n246), .A2(new_n248), .A3(new_n212), .A4(G68), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n281), .B2(new_n476), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n360), .A2(new_n361), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n557), .A2(new_n284), .B1(new_n364), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n546), .A2(new_n549), .A3(new_n550), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n284), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n360), .A2(new_n562), .A3(new_n361), .ZN(new_n563));
  AND2_X1   g0363(.A1(KEYINPUT15), .A2(G87), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT15), .A2(G87), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT77), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(new_n289), .A3(new_n292), .A4(new_n478), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n364), .A2(new_n558), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n561), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n543), .A2(new_n370), .A3(new_n469), .A4(new_n545), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n298), .B1(new_n547), .B2(new_n548), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n479), .A2(new_n348), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n364), .A2(new_n348), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT25), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n364), .A2(KEYINPUT81), .A3(KEYINPUT25), .A4(new_n348), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n575), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n250), .A2(new_n251), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n212), .A2(G87), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n212), .A2(G107), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT23), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n584), .A2(new_n434), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n540), .B1(new_n385), .B2(new_n590), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n591), .A2(G20), .ZN(new_n592));
  XNOR2_X1  g0392(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n587), .A2(new_n589), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT22), .B1(new_n349), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n589), .B1(new_n591), .B2(G20), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n599), .A3(new_n284), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G294), .ZN(new_n601));
  INV_X1    g0401(.A(G250), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n253), .ZN(new_n603));
  INV_X1    g0403(.A(G257), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n601), .B1(new_n392), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n259), .ZN(new_n608));
  OAI211_X1 g0408(.A(G264), .B(new_n258), .C1(new_n470), .C2(new_n544), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n508), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(G190), .A3(new_n508), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n583), .A2(new_n600), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n583), .A2(new_n600), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n298), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G179), .B2(new_n612), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n574), .B(new_n615), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n536), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n445), .A2(new_n499), .A3(new_n620), .ZN(G372));
  AND4_X1   g0421(.A1(new_n495), .A2(new_n497), .A3(new_n574), .A4(new_n615), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT78), .B1(new_n528), .B2(new_n501), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT21), .B1(new_n528), .B2(KEYINPUT78), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n531), .B2(new_n530), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n529), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n616), .A2(new_n618), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n573), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n485), .A2(new_n284), .ZN(new_n630));
  INV_X1    g0430(.A(new_n480), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n474), .A2(new_n298), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n574), .A2(new_n632), .A3(new_n633), .A4(new_n489), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n494), .A2(KEYINPUT26), .A3(new_n489), .A4(new_n574), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT82), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n640), .B(new_n629), .C1(new_n636), .C2(new_n637), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n628), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n445), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n426), .A2(new_n412), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n303), .A2(new_n304), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n369), .A2(new_n371), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n296), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n441), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n376), .B1(new_n650), .B2(new_n346), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(new_n651), .ZN(G369));
  AND2_X1   g0452(.A1(new_n212), .A2(G13), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n326), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n531), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n626), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n536), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT83), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT83), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT84), .ZN(new_n670));
  INV_X1    g0470(.A(new_n659), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n616), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n615), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n616), .A2(new_n670), .A3(new_n671), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(new_n627), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n627), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n669), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n675), .A2(new_n627), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n626), .A2(new_n671), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT85), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n680), .A2(new_n685), .A3(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n208), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n553), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n215), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n659), .B1(new_n628), .B2(new_n638), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n638), .B(KEYINPUT82), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n659), .B1(new_n697), .B2(new_n628), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n698), .B2(KEYINPUT29), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n454), .A2(new_n473), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G238), .A2(G1698), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n447), .B2(G1698), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n540), .B1(new_n702), .B2(new_n385), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n469), .B(new_n545), .C1(new_n703), .C2(new_n258), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n610), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n700), .A2(new_n530), .A3(KEYINPUT30), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n468), .A2(new_n471), .B1(new_n472), .B2(G270), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(new_n708), .A3(G179), .A4(new_n507), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n707), .B1(new_n709), .B2(new_n474), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n704), .A2(new_n370), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n474), .A2(new_n510), .A3(new_n612), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n713), .B2(new_n659), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n712), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT86), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT86), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(new_n717), .A3(new_n712), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n706), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n671), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n714), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT87), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n620), .A2(new_n499), .A3(new_n671), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n699), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n694), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n263), .B1(new_n653), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n689), .ZN(new_n734));
  AOI21_X1  g0534(.A(G330), .B1(new_n665), .B2(new_n666), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n669), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n662), .A2(new_n663), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n734), .B(KEYINPUT88), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n211), .B1(G20), .B2(new_n298), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n208), .A2(new_n385), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G45), .B2(new_n215), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n242), .B2(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n349), .A2(new_n207), .ZN(new_n748));
  INV_X1    g0548(.A(G355), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(G116), .B2(new_n207), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n744), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n212), .A2(new_n370), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n534), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n212), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n202), .B1(new_n434), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(G190), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n585), .B(new_n759), .C1(G68), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n534), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n212), .B1(new_n762), .B2(new_n370), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(KEYINPUT91), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(KEYINPUT91), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n757), .A2(new_n534), .A3(G200), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT90), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n761), .B1(new_n476), .B2(new_n767), .C1(new_n348), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n757), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n753), .A2(KEYINPUT89), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n753), .A2(KEYINPUT89), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(new_n762), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(new_n779), .A3(new_n773), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n777), .B1(new_n395), .B2(new_n780), .C1(new_n280), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n774), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n349), .B1(G329), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(new_n781), .C1(new_n786), .C2(new_n780), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G326), .A2(new_n755), .B1(new_n760), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n758), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n764), .A2(G294), .B1(new_n790), .B2(G303), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n789), .B(new_n791), .C1(new_n792), .C2(new_n771), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n772), .A2(new_n782), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n752), .B1(new_n794), .B2(new_n743), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n736), .B1(new_n740), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n366), .A2(new_n368), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n365), .B2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n646), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n369), .A2(new_n371), .A3(new_n671), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n698), .B(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n804), .A2(new_n728), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n728), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n734), .B(new_n805), .C1(KEYINPUT94), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT94), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n743), .A2(new_n737), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n742), .B1(G77), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G283), .A2(new_n760), .B1(new_n755), .B2(G303), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n348), .B2(new_n758), .ZN(new_n813));
  INV_X1    g0613(.A(new_n767), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G97), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n585), .B1(new_n785), .B2(new_n774), .C1(new_n780), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n781), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G116), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n771), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G87), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n815), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G137), .A2(new_n755), .B1(new_n760), .B2(G150), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT92), .B(G143), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n775), .B2(new_n781), .C1(new_n780), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n385), .B1(new_n774), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G58), .B2(new_n764), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n202), .B2(new_n758), .C1(new_n771), .C2(new_n288), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT93), .Z(new_n831));
  OAI21_X1  g0631(.A(new_n822), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n811), .B1(new_n832), .B2(new_n743), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n803), .B2(new_n738), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n808), .A2(new_n834), .ZN(G384));
  OAI211_X1 g0635(.A(G116), .B(new_n213), .C1(new_n483), .C2(KEYINPUT35), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(KEYINPUT35), .B2(new_n483), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT36), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n396), .A2(new_n215), .A3(new_n280), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n202), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(G13), .B(new_n326), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n713), .A2(new_n659), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT97), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n713), .A2(new_n845), .A3(new_n659), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n720), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT98), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT31), .B1(new_n843), .B2(KEYINPUT97), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(KEYINPUT98), .A3(new_n846), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n726), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n305), .B1(new_n295), .B2(new_n671), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n303), .A2(new_n304), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n659), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n802), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(KEYINPUT40), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n394), .A2(new_n400), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n403), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n420), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n409), .ZN(new_n862));
  INV_X1    g0662(.A(new_n657), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n442), .A2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n411), .B(new_n438), .C1(new_n415), .C2(new_n420), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n425), .A2(new_n657), .B1(new_n861), .B2(new_n409), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n389), .A2(new_n863), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n440), .B(new_n870), .C1(new_n421), .C2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT95), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n866), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n422), .A2(new_n863), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n441), .B2(new_n644), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n440), .B1(new_n421), .B2(new_n871), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n870), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n877), .A2(KEYINPUT100), .A3(new_n883), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n858), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT99), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n726), .A2(new_n852), .ZN(new_n890));
  INV_X1    g0690(.A(new_n846), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n845), .B1(new_n713), .B2(new_n659), .ZN(new_n892));
  NOR4_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(new_n848), .A4(KEYINPUT31), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT98), .B1(new_n850), .B2(new_n846), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n295), .A2(new_n671), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n855), .A2(new_n296), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n645), .A2(new_n671), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n803), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n889), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n866), .A2(new_n876), .A3(KEYINPUT96), .A4(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n869), .A2(new_n872), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT95), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n864), .B1(new_n427), .B2(new_n441), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n878), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT96), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n877), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n853), .A2(KEYINPUT99), .A3(new_n857), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n900), .A2(new_n901), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n888), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n445), .A3(new_n853), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  INV_X1    g0715(.A(new_n888), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n445), .A2(G330), .A3(new_n853), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n914), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n445), .B(new_n696), .C1(new_n698), .C2(KEYINPUT29), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n651), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n921), .B(new_n923), .Z(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n877), .A2(new_n925), .A3(new_n883), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n909), .A2(new_n901), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n925), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n645), .A2(new_n659), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n642), .A2(new_n671), .A3(new_n803), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n801), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n854), .A2(new_n856), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n927), .B1(new_n644), .B2(new_n863), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n326), .B2(new_n653), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n924), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n842), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n495), .A2(new_n497), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n632), .A2(new_n659), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n678), .A2(new_n682), .A3(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(KEYINPUT42), .B1(new_n492), .B2(new_n671), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(KEYINPUT42), .B2(new_n677), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n683), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n559), .A2(new_n550), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n659), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n574), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n629), .A2(new_n949), .A3(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT101), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n946), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n492), .A2(new_n659), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n944), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n680), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  INV_X1    g0764(.A(new_n957), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n946), .A2(new_n964), .A3(new_n965), .A4(new_n948), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n959), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT102), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT102), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n959), .A2(new_n969), .A3(new_n963), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n959), .A2(new_n966), .ZN(new_n971));
  INV_X1    g0771(.A(new_n963), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n689), .B(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n683), .A2(new_n684), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n962), .B1(new_n977), .B2(new_n686), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n687), .A2(new_n685), .A3(new_n961), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n687), .A2(KEYINPUT45), .A3(new_n685), .A4(new_n961), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n680), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n682), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n678), .B(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n665), .A2(KEYINPUT104), .A3(G330), .A4(new_n666), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n669), .A2(KEYINPUT104), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n990), .A2(new_n991), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT105), .A3(new_n730), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n980), .A2(new_n680), .A3(new_n985), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT105), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n995), .B1(new_n992), .B2(new_n993), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n729), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n988), .A2(new_n998), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n976), .B1(new_n1003), .B2(new_n730), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n974), .B1(new_n1004), .B2(new_n733), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n745), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n235), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n744), .B1(new_n207), .B2(new_n558), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n742), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n767), .A2(new_n288), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G77), .B2(new_n820), .ZN(new_n1011));
  INV_X1    g0811(.A(G137), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n349), .B1(new_n1012), .B2(new_n774), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n756), .A2(new_n824), .B1(new_n395), .B2(new_n758), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n780), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1014), .C1(G150), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n760), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n202), .A2(new_n781), .B1(new_n1017), .B2(new_n775), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT106), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n392), .B1(new_n774), .B2(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n756), .A2(new_n785), .B1(new_n348), .B2(new_n763), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G294), .C2(new_n760), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G283), .A2(new_n818), .B1(new_n1015), .B2(G303), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n790), .A2(G116), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT46), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n820), .A2(G97), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT47), .B1(new_n1020), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n743), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1020), .A2(new_n1029), .A3(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1009), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n739), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n957), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1005), .A2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n997), .A2(new_n730), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1001), .A2(new_n729), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n689), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n464), .B1(new_n288), .B2(new_n280), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n691), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT107), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n321), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT50), .B1(new_n321), .B2(new_n202), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n745), .B(new_n1047), .C1(new_n232), .C2(new_n464), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(G107), .B2(new_n207), .C1(new_n691), .C2(new_n748), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n741), .B1(new_n1049), .B2(new_n744), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n567), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n767), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n1028), .ZN(new_n1054));
  INV_X1    g0854(.A(G150), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n385), .B1(new_n774), .B2(new_n1055), .C1(new_n1017), .C2(new_n331), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n790), .A2(G77), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n756), .B2(new_n775), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n202), .A2(new_n780), .B1(new_n781), .B2(new_n288), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G311), .A2(new_n760), .B1(new_n755), .B2(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n502), .B2(new_n781), .C1(new_n1021), .C2(new_n780), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT48), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n792), .B2(new_n763), .C1(new_n816), .C2(new_n758), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n385), .B1(new_n783), .B2(G326), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n771), .B2(new_n512), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1060), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1050), .B1(new_n1031), .B2(new_n1070), .C1(new_n679), .C2(new_n1035), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1040), .B(new_n1071), .C1(new_n732), .C2(new_n1001), .ZN(G393));
  NAND2_X1  g0872(.A1(new_n962), .A2(new_n739), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n239), .A2(new_n1006), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n744), .B1(new_n476), .B2(new_n207), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n742), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n814), .A2(G77), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n818), .A2(new_n321), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n385), .B1(new_n774), .B2(new_n824), .C1(new_n288), .C2(new_n758), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G50), .B2(new_n760), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n821), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n775), .A2(new_n780), .B1(new_n756), .B2(new_n1055), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1015), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n585), .B1(new_n786), .B2(new_n774), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G294), .B2(new_n818), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n763), .A2(new_n512), .B1(new_n758), .B2(new_n792), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G303), .B2(new_n760), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(new_n348), .C2(new_n771), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1081), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1076), .B1(new_n1092), .B2(new_n743), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n988), .A2(new_n999), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n732), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT109), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n690), .B1(new_n1095), .B2(new_n1038), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n1003), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n980), .A2(new_n680), .A3(new_n985), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n680), .B1(new_n980), .B2(new_n985), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1038), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AND4_X1   g0903(.A1(new_n1098), .A2(new_n1003), .A3(new_n689), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1097), .B1(new_n1100), .B2(new_n1104), .ZN(G390));
  AND2_X1   g0905(.A1(new_n886), .A2(new_n887), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n929), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n801), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n695), .B2(new_n800), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n897), .A2(new_n898), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n727), .A2(G330), .A3(new_n803), .A4(new_n933), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n931), .B2(new_n801), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT110), .B1(new_n1114), .B2(new_n929), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n926), .C1(new_n925), .C2(new_n927), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1112), .B(new_n1113), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT110), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n934), .B2(new_n1107), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n928), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1119), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n853), .A2(G330), .A3(new_n857), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n732), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n742), .B1(new_n321), .B2(new_n810), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n928), .A2(new_n738), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n755), .A2(G283), .B1(new_n790), .B2(G87), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n348), .B2(new_n1017), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n585), .B1(new_n816), .B2(new_n774), .C1(new_n781), .C2(new_n476), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(G68), .C2(new_n820), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1077), .B1(new_n512), .B2(new_n780), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT112), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(KEYINPUT113), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1017), .A2(new_n1012), .B1(new_n756), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n585), .B(new_n1141), .C1(G125), .C2(new_n783), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n790), .A2(G150), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1143), .A2(KEYINPUT53), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n780), .A2(new_n827), .B1(new_n1143), .B2(KEYINPUT53), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT54), .B(G143), .Z(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1145), .C1(new_n818), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n820), .A2(G50), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n814), .A2(G159), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1142), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1138), .A2(KEYINPUT113), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1128), .B(new_n1129), .C1(new_n743), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1112), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1125), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n726), .B1(new_n722), .B2(new_n723), .ZN(new_n1158));
  AOI211_X1 g0958(.A(KEYINPUT87), .B(new_n714), .C1(new_n719), .C2(new_n721), .ZN(new_n1159));
  OAI211_X1 g0959(.A(G330), .B(new_n803), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1110), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1125), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n932), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n853), .A2(G330), .A3(new_n803), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1110), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1113), .A3(new_n1109), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n922), .A2(new_n651), .A3(new_n919), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT111), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT111), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n1168), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1157), .B(new_n1118), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1126), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1175), .A3(new_n689), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1154), .A2(new_n1176), .ZN(G378));
  OAI21_X1  g0977(.A(new_n1169), .B1(new_n1126), .B2(new_n1174), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n930), .A2(new_n935), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n863), .A2(new_n374), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n379), .B(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  AND4_X1   g0984(.A1(G330), .A2(new_n915), .A3(new_n916), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n913), .B2(G330), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n917), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n913), .A2(G330), .A3(new_n1184), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n936), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1178), .A2(KEYINPUT57), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT119), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT119), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1178), .A2(new_n1192), .A3(new_n1195), .A4(KEYINPUT57), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n689), .A3(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1187), .A2(KEYINPUT118), .A3(new_n1191), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT118), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1178), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n734), .B1(G50), .B2(new_n810), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1010), .B1(G116), .B2(new_n755), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT115), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n820), .A2(G58), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT114), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n385), .A2(G41), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1057), .B(new_n1208), .C1(new_n792), .C2(new_n774), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1051), .A2(new_n781), .B1(new_n780), .B2(new_n348), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G97), .C2(new_n760), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT58), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G33), .A2(G41), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1208), .A2(G50), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n755), .A2(G125), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1017), .B2(new_n827), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n790), .B2(new_n1146), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G128), .A2(new_n1015), .B1(new_n818), .B2(G137), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n1055), .C2(new_n767), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n783), .A2(G124), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1214), .B(new_n1223), .C1(new_n771), .C2(new_n775), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1215), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1213), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1203), .B1(new_n1227), .B2(new_n743), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1184), .B2(new_n738), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT117), .Z(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1200), .B2(new_n733), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1202), .A2(new_n1231), .ZN(G375));
  NOR2_X1   g1032(.A1(new_n781), .A2(new_n1055), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n385), .B1(new_n774), .B2(new_n1140), .C1(new_n775), .C2(new_n758), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n814), .C2(G50), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1207), .A2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT120), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G132), .A2(new_n755), .B1(new_n760), .B2(new_n1146), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1012), .B2(new_n780), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n585), .B1(new_n502), .B2(new_n774), .C1(new_n780), .C2(new_n792), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n756), .A2(new_n816), .B1(new_n476), .B2(new_n758), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G116), .B2(new_n760), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1053), .B(new_n1243), .C1(new_n280), .C2(new_n771), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1241), .B(new_n1244), .C1(G107), .C2(new_n818), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n743), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n741), .B1(new_n288), .B2(new_n809), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(new_n933), .C2(new_n738), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1167), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n732), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1168), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1174), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1253), .B2(new_n976), .ZN(G381));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G378), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1154), .A2(new_n1176), .A3(KEYINPUT121), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G375), .A2(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(G384), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1262), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n658), .A2(G213), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT122), .Z(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1260), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(new_n1268), .A3(G213), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT123), .ZN(G409));
  NAND3_X1  g1070(.A1(G390), .A2(new_n1036), .A3(new_n1005), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1099), .A2(new_n1098), .A3(new_n1003), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1003), .A2(new_n1103), .A3(new_n689), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT109), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1096), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1261), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1271), .A2(new_n1276), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1261), .A2(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(G387), .A3(new_n1275), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(G387), .B2(new_n1275), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(G390), .A2(KEYINPUT125), .A3(new_n1036), .A4(new_n1005), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1265), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1231), .C1(new_n1197), .C2(new_n1201), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1192), .A2(new_n733), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT118), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1192), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1187), .A2(new_n1191), .A3(KEYINPUT118), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1178), .A3(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1229), .B(new_n1292), .C1(new_n1296), .C2(new_n976), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1258), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1290), .B1(new_n1299), .B2(KEYINPUT124), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1253), .A2(KEYINPUT60), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1252), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n689), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1251), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n834), .A3(new_n808), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(G384), .A3(new_n1251), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1291), .A2(new_n1298), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1300), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1299), .A2(new_n1266), .A3(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  INV_X1    g1116(.A(G2897), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1266), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1265), .A2(new_n1317), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1319), .B1(new_n1308), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1267), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1315), .B(new_n1316), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1289), .B1(new_n1313), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1314), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1316), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1299), .A2(KEYINPUT124), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n1265), .A3(new_n1311), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1321), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1325), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1330), .A2(new_n1308), .ZN(new_n1333));
  OAI211_X1 g1133(.A(KEYINPUT127), .B(new_n1328), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1321), .B1(new_n1300), .B2(new_n1311), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1312), .B1(new_n1336), .B2(new_n1325), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT127), .B1(new_n1337), .B2(new_n1328), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1324), .B1(new_n1335), .B2(new_n1338), .ZN(G405));
  AOI21_X1  g1139(.A(new_n1259), .B1(new_n1202), .B2(new_n1231), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1291), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1308), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1289), .ZN(G402));
endmodule


