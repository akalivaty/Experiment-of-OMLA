//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT64), .B2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n458), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n458), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n465), .B2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n458), .A2(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n474), .A2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n459), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n458), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n485), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n489), .B1(new_n475), .B2(new_n476), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n460), .A2(new_n461), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n487), .A2(new_n501), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n495), .A2(new_n496), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n479), .B2(G126), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT65), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n516), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT66), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n512), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n524), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n515), .A2(G51), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT67), .B(G89), .Z(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n519), .A2(new_n520), .B1(new_n513), .B2(new_n514), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(G90), .B1(new_n515), .B2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT68), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n540), .A2(new_n547), .A3(KEYINPUT68), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n512), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n515), .A2(G43), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT69), .B(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n523), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT70), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  AND2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n522), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n519), .B2(new_n520), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n521), .A2(new_n522), .A3(G91), .ZN(new_n577));
  AND4_X1   g152(.A1(new_n564), .A2(new_n571), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G65), .B1(new_n542), .B2(new_n543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(new_n574), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n539), .B2(G91), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n564), .B1(new_n581), .B2(new_n571), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  OR2_X1    g159(.A1(new_n533), .A2(new_n537), .ZN(G286));
  NAND2_X1  g160(.A1(new_n539), .A2(G87), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT72), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n521), .A2(G74), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n515), .B2(G49), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n515), .A2(G48), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT73), .B1(new_n544), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n521), .A2(new_n596), .A3(G61), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n593), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n539), .A2(G86), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT74), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n521), .A2(new_n522), .A3(G86), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT74), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n539), .A2(G85), .B1(new_n515), .B2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n512), .B2(new_n609), .ZN(G290));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n523), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n544), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n618), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(G301), .B(new_n622), .S(new_n623), .Z(G284));
  MUX2_X1   g199(.A(G301), .B(new_n622), .S(new_n623), .Z(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(new_n622), .ZN(new_n630));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G860), .ZN(G148));
  OAI21_X1  g207(.A(new_n623), .B1(new_n553), .B2(new_n556), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n622), .A2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n492), .A2(new_n469), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT76), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n477), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n479), .A2(G123), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n644), .A2(new_n458), .A3(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n458), .B2(G111), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G2104), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n642), .B(new_n643), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n641), .A2(new_n650), .A3(new_n651), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(KEYINPUT79), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n673), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n670), .B1(new_n672), .B2(new_n673), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n670), .A2(new_n671), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n687), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n687), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT80), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G33), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT25), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n477), .A2(G139), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT85), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n492), .A2(G127), .ZN(new_n712));
  AND2_X1   g287(.A1(G115), .A2(G2104), .ZN(new_n713));
  OAI21_X1  g288(.A(G2105), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT86), .Z(new_n716));
  OAI21_X1  g291(.A(new_n706), .B1(new_n716), .B2(new_n705), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2072), .Z(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G105), .B2(new_n469), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n477), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT88), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G29), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT81), .B(G29), .Z(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G34), .B2(new_n732), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G160), .B2(G29), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n729), .A2(new_n730), .B1(G2084), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n718), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n731), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT84), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G116), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT83), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n477), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n479), .A2(G128), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n742), .B1(G29), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2067), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT30), .B(G28), .Z(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G29), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n649), .A2(new_n731), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(new_n755), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT91), .Z(new_n759));
  INV_X1    g334(.A(new_n731), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G27), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n760), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2078), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n557), .B2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G21), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G168), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n770), .C1(G2084), .C2(new_n735), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n751), .A2(new_n759), .A3(new_n763), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n760), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n760), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  INV_X1    g354(.A(G16), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G4), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n622), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1348), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n627), .B2(new_n780), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n782), .A2(new_n783), .B1(new_n786), .B2(G1956), .ZN(new_n787));
  NOR2_X1   g362(.A1(G5), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G171), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n776), .A2(new_n777), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n730), .B2(new_n729), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n782), .A2(new_n783), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n786), .A2(G1956), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n792), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n772), .A2(new_n779), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n718), .A2(KEYINPUT89), .A3(new_n736), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n739), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n739), .A2(new_n798), .A3(new_n802), .A4(new_n799), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(new_n780), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n780), .B2(G23), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n780), .A2(G22), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n780), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1971), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(G6), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G305), .B2(new_n780), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n816), .A2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT34), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n814), .A2(new_n823), .A3(new_n819), .A4(new_n820), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G24), .ZN(new_n825));
  XOR2_X1   g400(.A(G290), .B(KEYINPUT82), .Z(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1986), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n477), .A2(G131), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n479), .A2(G119), .ZN(new_n830));
  OR2_X1    g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  MUX2_X1   g408(.A(G25), .B(new_n833), .S(new_n760), .Z(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n822), .A2(new_n824), .A3(new_n828), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n801), .A2(new_n803), .B1(new_n838), .B2(new_n839), .ZN(G311));
  NAND2_X1  g415(.A1(new_n801), .A2(new_n803), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(G150));
  NOR2_X1   g418(.A1(new_n622), .A2(new_n631), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n512), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n515), .A2(G55), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT95), .B(G93), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n523), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n557), .A2(new_n851), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n556), .A2(new_n553), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n845), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(G860), .B1(new_n847), .B2(new_n850), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n504), .A2(new_n506), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n749), .B(new_n863), .Z(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n749), .B(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT97), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n726), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n715), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n726), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n727), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n716), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n638), .B(new_n833), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n477), .A2(G142), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT98), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n479), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n458), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n879), .B(new_n885), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n876), .A2(new_n878), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n872), .A2(new_n877), .A3(new_n874), .A4(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(G160), .B(KEYINPUT96), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n649), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n878), .A2(new_n887), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n877), .B1(new_n872), .B2(new_n874), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n893), .B(new_n889), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n896), .A4(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n896), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n893), .B1(new_n888), .B2(new_n889), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n900), .A2(new_n904), .ZN(G395));
  XNOR2_X1  g480(.A(new_n634), .B(new_n855), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n578), .B2(new_n582), .ZN(new_n907));
  INV_X1    g482(.A(new_n620), .ZN(new_n908));
  INV_X1    g483(.A(new_n571), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n576), .A2(new_n577), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT71), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n581), .A2(new_n564), .A3(new_n571), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n908), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(G299), .A2(new_n912), .A3(new_n620), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n915), .B2(new_n916), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT101), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n918), .B1(new_n926), .B2(new_n906), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(G288), .B(G305), .ZN(new_n929));
  XNOR2_X1  g504(.A(G303), .B(G290), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n929), .B(new_n930), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n928), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g511(.A(new_n935), .B1(G868), .B2(new_n851), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(new_n550), .ZN(new_n940));
  OAI21_X1  g515(.A(G168), .B1(new_n940), .B2(new_n548), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n549), .A2(G286), .A3(new_n550), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n855), .A2(KEYINPUT103), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n854), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(KEYINPUT102), .A3(new_n854), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT102), .B1(new_n945), .B2(new_n854), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n943), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n917), .A2(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n925), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n945), .B(new_n855), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n916), .A3(new_n915), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT104), .B(new_n950), .C1(new_n953), .C2(new_n954), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n961), .B2(new_n931), .ZN(new_n962));
  INV_X1    g537(.A(new_n931), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n957), .A2(new_n963), .A3(new_n959), .A4(new_n960), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n939), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n959), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT104), .B1(new_n926), .B2(new_n950), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n966), .A2(new_n967), .A3(new_n931), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n950), .A2(new_n917), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n958), .B1(new_n952), .B2(new_n951), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n931), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n896), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n968), .A2(KEYINPUT43), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n938), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n966), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT43), .B1(new_n976), .B2(new_n963), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n938), .B1(new_n977), .B2(new_n962), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n968), .B2(new_n972), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n931), .B1(new_n966), .B2(new_n967), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(new_n964), .A3(new_n939), .A4(new_n896), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n975), .A2(new_n979), .A3(KEYINPUT44), .A4(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n493), .B2(new_n498), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G125), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n491), .B2(new_n459), .ZN(new_n990));
  INV_X1    g565(.A(new_n463), .ZN(new_n991));
  OAI21_X1  g566(.A(G2105), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(G40), .A3(new_n467), .A4(new_n470), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n749), .B(G2067), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n998), .B2(new_n726), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n994), .A2(G1996), .A3(new_n726), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT106), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n727), .A2(new_n995), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n994), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n833), .B(new_n835), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(KEYINPUT107), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(KEYINPUT107), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n994), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n994), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT48), .Z(new_n1014));
  OAI21_X1  g589(.A(new_n1001), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n835), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n833), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT126), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G2067), .B2(new_n749), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n994), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT127), .Z(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n568), .B2(new_n570), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n910), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n568), .A2(new_n570), .A3(new_n1025), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n581), .A2(KEYINPUT57), .A3(new_n571), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1026), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n581), .A3(new_n1028), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1023), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1030), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G40), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n464), .A2(new_n471), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n504), .B2(new_n506), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n499), .B2(new_n507), .ZN(new_n1044));
  AOI22_X1  g619(.A1(KEYINPUT111), .A2(new_n1043), .B1(new_n1044), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1956), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n993), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(G2072), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1051), .C1(new_n1044), .C2(KEYINPUT45), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1038), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1038), .B(KEYINPUT117), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1040), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n508), .A2(new_n985), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(KEYINPUT50), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1061));
  OAI22_X1  g636(.A1(new_n1060), .A2(G1348), .B1(G2067), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n908), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1044), .A2(new_n1042), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1047), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1052), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1054), .A2(new_n1073), .A3(new_n1071), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1054), .B2(new_n1073), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1061), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1061), .A2(KEYINPUT119), .A3(new_n1077), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1049), .B(new_n995), .C1(new_n1044), .C2(KEYINPUT45), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1080), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n557), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g663(.A(new_n908), .B1(G2067), .B2(new_n1061), .C1(new_n1060), .C2(G1348), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT120), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n557), .B(new_n1092), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1062), .A2(new_n620), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n1089), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1088), .A2(new_n1090), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1072), .B1(new_n1076), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G303), .A2(G8), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT55), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1058), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n777), .C1(new_n1044), .C2(new_n1042), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1049), .B1(new_n1044), .B2(KEYINPUT45), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT108), .ZN(new_n1105));
  INV_X1    g680(.A(G1971), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT108), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1049), .B(new_n1107), .C1(new_n1044), .C2(KEYINPUT45), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1103), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1105), .A2(KEYINPUT109), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1098), .B(new_n1100), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1098), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(G288), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT52), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n804), .B2(G1976), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(new_n1116), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT110), .ZN(new_n1121));
  INV_X1    g696(.A(G1981), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n600), .A2(new_n606), .A3(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n603), .B(new_n593), .C1(new_n599), .C2(G651), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1123), .B(KEYINPUT49), .C1(new_n1124), .C2(new_n1122), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1114), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(new_n600), .B2(new_n601), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT49), .B1(new_n1128), .B2(new_n1123), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1121), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT49), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1123), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1127), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(KEYINPUT110), .A3(new_n1114), .A4(new_n1125), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1120), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1100), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1045), .A2(new_n777), .A3(new_n1047), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1098), .B1(new_n1109), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n1140));
  NAND3_X1  g715(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(G168), .B2(new_n1098), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1144), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT112), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT45), .B1(new_n863), .B2(new_n985), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n993), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT112), .B(new_n1040), .C1(new_n1041), .C2(KEYINPUT45), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n493), .A2(new_n498), .A3(new_n485), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT65), .B1(new_n504), .B2(new_n506), .ZN(new_n1154));
  OAI211_X1 g729(.A(KEYINPUT45), .B(new_n985), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G2084), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1156), .A2(new_n769), .B1(new_n1060), .B2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1147), .B(new_n1148), .C1(new_n1158), .C2(new_n1098), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1152), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT112), .B1(new_n988), .B2(new_n1040), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n769), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1060), .A2(new_n1157), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1144), .B1(new_n1164), .B2(G8), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1146), .B1(new_n1158), .B2(new_n1148), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1113), .A2(new_n1139), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1169));
  INV_X1    g744(.A(G2078), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1060), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1171), .A2(new_n1172), .B1(new_n790), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(KEYINPUT53), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n1040), .A3(new_n988), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1174), .A2(new_n1175), .A3(G301), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1156), .A2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1173), .A2(new_n790), .ZN(new_n1182));
  AOI21_X1  g757(.A(G2078), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1181), .B(new_n1182), .C1(new_n1183), .C2(KEYINPUT53), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(G171), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1182), .B(new_n1178), .C1(new_n1183), .C2(KEYINPUT53), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT123), .B1(new_n1187), .B2(G171), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1179), .B(new_n1180), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1180), .B1(new_n1187), .B2(G171), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(G171), .B2(new_n1184), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1097), .A2(new_n1168), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1164), .A2(new_n1193), .A3(G8), .A4(G168), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1109), .A2(new_n1137), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(G8), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1194), .B1(new_n1196), .B2(new_n1100), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1135), .B1(new_n1113), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1199), .A2(new_n1112), .A3(new_n1102), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1136), .B1(new_n1200), .B2(G8), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1158), .A2(new_n1098), .A3(G286), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1135), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT63), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g779(.A(G1976), .B(G288), .C1(new_n1130), .C2(new_n1134), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1114), .B1(new_n1205), .B2(new_n1132), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1198), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1167), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1208), .A2(new_n1209), .A3(KEYINPUT62), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1113), .A2(new_n1139), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n1212));
  OAI21_X1  g787(.A(KEYINPUT124), .B1(new_n1167), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1185), .B1(new_n1167), .B2(new_n1212), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1192), .A2(new_n1207), .A3(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g791(.A(G290), .B(G1986), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1011), .B1(new_n994), .B2(new_n1217), .ZN(new_n1218));
  AND3_X1   g793(.A1(new_n1216), .A2(KEYINPUT125), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(KEYINPUT125), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1022), .B1(new_n1219), .B2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g796(.A1(new_n684), .A2(G319), .ZN(new_n1223));
  NOR3_X1   g797(.A1(G229), .A2(G401), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1224), .B1(new_n902), .B2(new_n903), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n965), .A2(new_n973), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  OR2_X1    g801(.A1(new_n1225), .A2(new_n1226), .ZN(G225));
endmodule


