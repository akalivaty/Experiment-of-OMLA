

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775;

  INV_X1 U368 ( .A(G953), .ZN(n762) );
  BUF_X2 U369 ( .A(n679), .Z(n687) );
  NOR2_X2 U370 ( .A1(n755), .A2(G953), .ZN(n756) );
  XNOR2_X2 U371 ( .A(n471), .B(n440), .ZN(n670) );
  XNOR2_X2 U372 ( .A(n438), .B(G128), .ZN(n482) );
  XNOR2_X2 U373 ( .A(G478), .B(n515), .ZN(n568) );
  XNOR2_X2 U374 ( .A(n462), .B(KEYINPUT75), .ZN(n554) );
  AND2_X2 U375 ( .A1(n725), .A2(n726), .ZN(n462) );
  NOR2_X1 U376 ( .A1(n627), .A2(n600), .ZN(n601) );
  NOR2_X1 U377 ( .A1(n416), .A2(n413), .ZN(n420) );
  XNOR2_X1 U378 ( .A(n365), .B(KEYINPUT106), .ZN(n596) );
  BUF_X1 U379 ( .A(n558), .Z(n559) );
  NOR2_X1 U380 ( .A1(n729), .A2(n728), .ZN(n726) );
  XNOR2_X1 U381 ( .A(n393), .B(n392), .ZN(n591) );
  XNOR2_X1 U382 ( .A(n461), .B(n460), .ZN(n729) );
  OR2_X1 U383 ( .A1(n649), .A2(n490), .ZN(n493) );
  XNOR2_X1 U384 ( .A(n370), .B(n452), .ZN(n681) );
  XNOR2_X1 U385 ( .A(n503), .B(n484), .ZN(n471) );
  INV_X1 U386 ( .A(KEYINPUT60), .ZN(n348) );
  INV_X1 U387 ( .A(KEYINPUT56), .ZN(n346) );
  INV_X1 U388 ( .A(G143), .ZN(n438) );
  XNOR2_X1 U389 ( .A(KEYINPUT68), .B(G101), .ZN(n464) );
  NAND2_X1 U390 ( .A1(n763), .A2(n672), .ZN(n345) );
  NAND2_X1 U391 ( .A1(n763), .A2(n672), .ZN(n746) );
  XNOR2_X1 U392 ( .A(n347), .B(n346), .ZN(G51) );
  NAND2_X1 U393 ( .A1(n652), .A2(n682), .ZN(n347) );
  XNOR2_X1 U394 ( .A(n349), .B(n348), .ZN(G60) );
  NAND2_X1 U395 ( .A1(n647), .A2(n682), .ZN(n349) );
  NOR2_X1 U396 ( .A1(n709), .A2(n625), .ZN(n366) );
  NAND2_X1 U397 ( .A1(n381), .A2(n382), .ZN(n380) );
  AND2_X1 U398 ( .A1(n654), .A2(n547), .ZN(n548) );
  NOR2_X1 U399 ( .A1(G237), .A2(G953), .ZN(n466) );
  XNOR2_X1 U400 ( .A(n376), .B(n375), .ZN(n478) );
  XNOR2_X1 U401 ( .A(G116), .B(G113), .ZN(n376) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(G119), .ZN(n375) );
  XNOR2_X1 U403 ( .A(n435), .B(n436), .ZN(n757) );
  XNOR2_X1 U404 ( .A(n434), .B(G110), .ZN(n436) );
  INV_X1 U405 ( .A(KEYINPUT93), .ZN(n434) );
  NOR2_X1 U406 ( .A1(n423), .A2(n418), .ZN(n417) );
  INV_X1 U407 ( .A(n426), .ZN(n418) );
  INV_X1 U408 ( .A(KEYINPUT38), .ZN(n369) );
  XNOR2_X1 U409 ( .A(n380), .B(n379), .ZN(n378) );
  XNOR2_X1 U410 ( .A(n366), .B(KEYINPUT70), .ZN(n383) );
  INV_X1 U411 ( .A(KEYINPUT46), .ZN(n379) );
  INV_X1 U412 ( .A(KEYINPUT48), .ZN(n377) );
  AND2_X1 U413 ( .A1(n672), .A2(n364), .ZN(n403) );
  NAND2_X1 U414 ( .A1(n359), .A2(n390), .ZN(n389) );
  NOR2_X1 U415 ( .A1(n613), .A2(KEYINPUT28), .ZN(n390) );
  NAND2_X1 U416 ( .A1(n613), .A2(KEYINPUT28), .ZN(n388) );
  XNOR2_X1 U417 ( .A(n441), .B(G469), .ZN(n558) );
  INV_X1 U418 ( .A(G902), .ZN(n497) );
  XNOR2_X1 U419 ( .A(n558), .B(KEYINPUT1), .ZN(n725) );
  XNOR2_X1 U420 ( .A(n471), .B(n472), .ZN(n664) );
  XOR2_X1 U421 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n447) );
  XNOR2_X1 U422 ( .A(G146), .B(KEYINPUT78), .ZN(n432) );
  XNOR2_X1 U423 ( .A(n351), .B(n431), .ZN(n396) );
  XNOR2_X1 U424 ( .A(n757), .B(n437), .ZN(n479) );
  OR2_X1 U425 ( .A1(n359), .A2(n391), .ZN(n387) );
  INV_X1 U426 ( .A(n591), .ZN(n731) );
  XNOR2_X1 U427 ( .A(n541), .B(n362), .ZN(n551) );
  XNOR2_X1 U428 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U429 ( .A1(G902), .A2(n681), .ZN(n461) );
  XNOR2_X1 U430 ( .A(n457), .B(n456), .ZN(n458) );
  BUF_X1 U431 ( .A(n725), .Z(n374) );
  INV_X1 U432 ( .A(n502), .ZN(n422) );
  NAND2_X1 U433 ( .A1(n502), .A2(n424), .ZN(n423) );
  NOR2_X1 U434 ( .A1(n495), .A2(KEYINPUT19), .ZN(n426) );
  NAND2_X1 U435 ( .A1(n429), .A2(KEYINPUT0), .ZN(n411) );
  NAND2_X1 U436 ( .A1(n415), .A2(n414), .ZN(n413) );
  AND2_X1 U437 ( .A1(n421), .A2(n355), .ZN(n414) );
  NAND2_X1 U438 ( .A1(n427), .A2(n417), .ZN(n415) );
  NAND2_X1 U439 ( .A1(n422), .A2(KEYINPUT0), .ZN(n421) );
  NOR2_X1 U440 ( .A1(n430), .A2(n423), .ZN(n416) );
  XNOR2_X1 U441 ( .A(G137), .B(G146), .ZN(n467) );
  XNOR2_X1 U442 ( .A(KEYINPUT5), .B(G131), .ZN(n463) );
  INV_X1 U443 ( .A(KEYINPUT90), .ZN(n573) );
  XNOR2_X1 U444 ( .A(G119), .B(G140), .ZN(n446) );
  XOR2_X1 U445 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n505) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT9), .ZN(n504) );
  XNOR2_X1 U447 ( .A(G116), .B(G107), .ZN(n507) );
  XNOR2_X1 U448 ( .A(n485), .B(KEYINPUT10), .ZN(n523) );
  NAND2_X1 U449 ( .A1(n714), .A2(n713), .ZN(n719) );
  INV_X1 U450 ( .A(n631), .ZN(n427) );
  INV_X1 U451 ( .A(n430), .ZN(n412) );
  INV_X1 U452 ( .A(G237), .ZN(n491) );
  XNOR2_X1 U453 ( .A(G902), .B(KEYINPUT15), .ZN(n638) );
  XNOR2_X1 U454 ( .A(n533), .B(n532), .ZN(n569) );
  XNOR2_X1 U455 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U456 ( .A1(G902), .A2(n643), .ZN(n533) );
  AND2_X1 U457 ( .A1(n634), .A2(n356), .ZN(n672) );
  XNOR2_X1 U458 ( .A(n368), .B(n377), .ZN(n634) );
  XNOR2_X1 U459 ( .A(n482), .B(n439), .ZN(n503) );
  INV_X1 U460 ( .A(G134), .ZN(n439) );
  XOR2_X1 U461 ( .A(G122), .B(G104), .Z(n525) );
  XNOR2_X1 U462 ( .A(G143), .B(G113), .ZN(n524) );
  XNOR2_X1 U463 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n517) );
  XNOR2_X1 U464 ( .A(n522), .B(n523), .ZN(n527) );
  XNOR2_X1 U465 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n484) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n476) );
  XNOR2_X1 U467 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n481) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U469 ( .A(n585), .B(KEYINPUT39), .ZN(n626) );
  AND2_X1 U470 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U471 ( .A(G472), .ZN(n392) );
  NAND2_X1 U472 ( .A1(n664), .A2(n497), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n451), .B(n454), .ZN(n370) );
  XNOR2_X1 U474 ( .A(G128), .B(G110), .ZN(n449) );
  XNOR2_X1 U475 ( .A(n670), .B(n394), .ZN(n689) );
  XNOR2_X1 U476 ( .A(n479), .B(n395), .ZN(n394) );
  XNOR2_X1 U477 ( .A(n396), .B(n433), .ZN(n395) );
  NOR2_X1 U478 ( .A1(n385), .A2(n384), .ZN(n605) );
  INV_X1 U479 ( .A(KEYINPUT36), .ZN(n367) );
  XNOR2_X1 U480 ( .A(n545), .B(KEYINPUT32), .ZN(n654) );
  OR2_X1 U481 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U482 ( .A(n607), .B(n606), .ZN(n701) );
  INV_X1 U483 ( .A(KEYINPUT82), .ZN(n606) );
  NAND2_X1 U484 ( .A1(n352), .A2(n386), .ZN(n607) );
  AND2_X1 U485 ( .A1(n387), .A2(n604), .ZN(n386) );
  AND2_X1 U486 ( .A1(n388), .A2(n559), .ZN(n350) );
  XNOR2_X1 U487 ( .A(G137), .B(KEYINPUT69), .ZN(n351) );
  AND2_X1 U488 ( .A1(n389), .A2(n350), .ZN(n352) );
  XOR2_X1 U489 ( .A(KEYINPUT79), .B(KEYINPUT94), .Z(n353) );
  OR2_X1 U490 ( .A1(n374), .A2(n546), .ZN(n354) );
  OR2_X1 U491 ( .A1(n423), .A2(n429), .ZN(n355) );
  AND2_X1 U492 ( .A1(n633), .A2(n662), .ZN(n356) );
  AND2_X1 U493 ( .A1(n401), .A2(n618), .ZN(n357) );
  OR2_X1 U494 ( .A1(n574), .A2(KEYINPUT44), .ZN(n358) );
  XOR2_X1 U495 ( .A(G131), .B(G140), .Z(n522) );
  NOR2_X1 U496 ( .A1(n594), .A2(n591), .ZN(n359) );
  NOR2_X1 U497 ( .A1(n551), .A2(n354), .ZN(n360) );
  OR2_X1 U498 ( .A1(n556), .A2(KEYINPUT34), .ZN(n361) );
  INV_X1 U499 ( .A(KEYINPUT28), .ZN(n391) );
  XOR2_X1 U500 ( .A(n540), .B(n539), .Z(n362) );
  NAND2_X1 U501 ( .A1(n637), .A2(n639), .ZN(n363) );
  NAND2_X1 U502 ( .A1(n635), .A2(n639), .ZN(n364) );
  NAND2_X1 U503 ( .A1(n569), .A2(n568), .ZN(n365) );
  XNOR2_X1 U504 ( .A(n601), .B(n367), .ZN(n602) );
  XNOR2_X1 U505 ( .A(n529), .B(n528), .ZN(n643) );
  NAND2_X1 U506 ( .A1(n378), .A2(n383), .ZN(n368) );
  XNOR2_X1 U507 ( .A(n631), .B(n369), .ZN(n588) );
  XNOR2_X2 U508 ( .A(n493), .B(n492), .ZN(n631) );
  XNOR2_X1 U509 ( .A(n589), .B(KEYINPUT41), .ZN(n749) );
  NAND2_X1 U510 ( .A1(n371), .A2(n361), .ZN(n400) );
  INV_X1 U511 ( .A(n750), .ZN(n371) );
  XNOR2_X2 U512 ( .A(n475), .B(KEYINPUT33), .ZN(n750) );
  NAND2_X1 U513 ( .A1(n397), .A2(n357), .ZN(n535) );
  NOR2_X2 U514 ( .A1(n554), .A2(n597), .ZN(n475) );
  XNOR2_X2 U515 ( .A(n372), .B(n640), .ZN(n679) );
  NAND2_X1 U516 ( .A1(n402), .A2(n404), .ZN(n372) );
  XNOR2_X1 U517 ( .A(n373), .B(n573), .ZN(n575) );
  NAND2_X1 U518 ( .A1(n571), .A2(n572), .ZN(n373) );
  NAND2_X1 U519 ( .A1(n660), .A2(n706), .ZN(n406) );
  INV_X1 U520 ( .A(n775), .ZN(n381) );
  INV_X1 U521 ( .A(n772), .ZN(n382) );
  INV_X1 U522 ( .A(n389), .ZN(n384) );
  NAND2_X1 U523 ( .A1(n387), .A2(n350), .ZN(n385) );
  NAND2_X1 U524 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U525 ( .A1(n750), .A2(n399), .ZN(n398) );
  INV_X1 U526 ( .A(KEYINPUT34), .ZN(n399) );
  NAND2_X1 U527 ( .A1(n556), .A2(KEYINPUT34), .ZN(n401) );
  NAND2_X1 U528 ( .A1(n345), .A2(n363), .ZN(n402) );
  NAND2_X1 U529 ( .A1(n403), .A2(n763), .ZN(n404) );
  XNOR2_X1 U530 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X2 U531 ( .A(n577), .B(n576), .ZN(n763) );
  NAND2_X1 U532 ( .A1(n655), .A2(n405), .ZN(n570) );
  NAND2_X1 U533 ( .A1(n406), .A2(n611), .ZN(n405) );
  XNOR2_X2 U534 ( .A(n565), .B(n564), .ZN(n660) );
  NAND2_X1 U535 ( .A1(n407), .A2(n553), .ZN(n655) );
  XNOR2_X1 U536 ( .A(n552), .B(n408), .ZN(n407) );
  INV_X1 U537 ( .A(KEYINPUT89), .ZN(n408) );
  NOR2_X1 U538 ( .A1(n412), .A2(n409), .ZN(n428) );
  INV_X1 U539 ( .A(n429), .ZN(n409) );
  NAND2_X1 U540 ( .A1(n410), .A2(n425), .ZN(n419) );
  NAND2_X1 U541 ( .A1(n427), .A2(n426), .ZN(n425) );
  NOR2_X1 U542 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U543 ( .A1(n428), .A2(n425), .ZN(n604) );
  NAND2_X1 U544 ( .A1(n420), .A2(n419), .ZN(n560) );
  INV_X1 U545 ( .A(KEYINPUT0), .ZN(n424) );
  NAND2_X1 U546 ( .A1(n427), .A2(n713), .ZN(n600) );
  NAND2_X1 U547 ( .A1(n495), .A2(KEYINPUT19), .ZN(n429) );
  NAND2_X1 U548 ( .A1(n631), .A2(KEYINPUT19), .ZN(n430) );
  XNOR2_X1 U549 ( .A(n523), .B(n351), .ZN(n671) );
  INV_X1 U550 ( .A(n522), .ZN(n440) );
  INV_X1 U551 ( .A(KEYINPUT47), .ZN(n608) );
  INV_X1 U552 ( .A(n360), .ZN(n547) );
  INV_X1 U553 ( .A(KEYINPUT24), .ZN(n445) );
  INV_X1 U554 ( .A(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U555 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U556 ( .A(n509), .B(n508), .ZN(n510) );
  BUF_X1 U557 ( .A(n560), .Z(n556) );
  NOR2_X1 U558 ( .A1(n603), .A2(n602), .ZN(n709) );
  NAND2_X1 U559 ( .A1(n762), .A2(G227), .ZN(n431) );
  XNOR2_X1 U560 ( .A(n353), .B(n432), .ZN(n433) );
  XNOR2_X1 U561 ( .A(G107), .B(G104), .ZN(n435) );
  XNOR2_X1 U562 ( .A(n464), .B(KEYINPUT72), .ZN(n437) );
  NAND2_X1 U563 ( .A1(n689), .A2(n497), .ZN(n441) );
  XOR2_X1 U564 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n443) );
  NAND2_X1 U565 ( .A1(G234), .A2(n638), .ZN(n442) );
  XNOR2_X1 U566 ( .A(n443), .B(n442), .ZN(n455) );
  NAND2_X1 U567 ( .A1(n455), .A2(G221), .ZN(n444) );
  XNOR2_X1 U568 ( .A(n444), .B(KEYINPUT21), .ZN(n728) );
  XNOR2_X1 U569 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U570 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X2 U572 ( .A(G146), .B(G125), .ZN(n485) );
  INV_X1 U573 ( .A(n671), .ZN(n451) );
  NAND2_X1 U574 ( .A1(n762), .A2(G234), .ZN(n453) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(n453), .Z(n512) );
  NAND2_X1 U576 ( .A1(G221), .A2(n512), .ZN(n454) );
  NAND2_X1 U577 ( .A1(G217), .A2(n455), .ZN(n459) );
  XOR2_X1 U578 ( .A(KEYINPUT96), .B(KEYINPUT77), .Z(n457) );
  XNOR2_X1 U579 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U580 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U581 ( .A(n478), .B(n465), .ZN(n470) );
  XNOR2_X1 U582 ( .A(n466), .B(KEYINPUT76), .ZN(n516) );
  NAND2_X1 U583 ( .A1(G210), .A2(n516), .ZN(n468) );
  XNOR2_X1 U584 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U585 ( .A(n470), .B(n469), .ZN(n472) );
  INV_X1 U586 ( .A(KEYINPUT107), .ZN(n473) );
  XNOR2_X1 U587 ( .A(n473), .B(KEYINPUT6), .ZN(n474) );
  XNOR2_X1 U588 ( .A(n731), .B(n474), .ZN(n597) );
  XNOR2_X1 U589 ( .A(n476), .B(KEYINPUT74), .ZN(n477) );
  XNOR2_X1 U590 ( .A(n478), .B(n477), .ZN(n759) );
  XNOR2_X1 U591 ( .A(n479), .B(n759), .ZN(n489) );
  NAND2_X1 U592 ( .A1(n762), .A2(G224), .ZN(n480) );
  XNOR2_X1 U593 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n482), .B(n483), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U597 ( .A(n489), .B(n488), .ZN(n649) );
  INV_X1 U598 ( .A(n638), .ZN(n490) );
  NAND2_X1 U599 ( .A1(n497), .A2(n491), .ZN(n494) );
  NAND2_X1 U600 ( .A1(n494), .A2(G210), .ZN(n492) );
  NAND2_X1 U601 ( .A1(n494), .A2(G214), .ZN(n713) );
  INV_X1 U602 ( .A(n713), .ZN(n495) );
  XNOR2_X1 U603 ( .A(KEYINPUT14), .B(n496), .ZN(n712) );
  NAND2_X1 U604 ( .A1(n497), .A2(G953), .ZN(n499) );
  OR2_X1 U605 ( .A1(G953), .A2(G952), .ZN(n498) );
  AND2_X1 U606 ( .A1(n499), .A2(n498), .ZN(n500) );
  AND2_X1 U607 ( .A1(n712), .A2(n500), .ZN(n579) );
  NAND2_X1 U608 ( .A1(G953), .A2(G898), .ZN(n501) );
  AND2_X1 U609 ( .A1(n579), .A2(n501), .ZN(n502) );
  INV_X1 U610 ( .A(n503), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n509) );
  XNOR2_X1 U612 ( .A(n511), .B(n510), .ZN(n514) );
  NAND2_X1 U613 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n514), .B(n513), .ZN(n684) );
  NOR2_X1 U615 ( .A1(G902), .A2(n684), .ZN(n515) );
  NAND2_X1 U616 ( .A1(n516), .A2(G214), .ZN(n520) );
  XOR2_X1 U617 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n518) );
  XNOR2_X1 U618 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U620 ( .A(n521), .B(KEYINPUT100), .Z(n529) );
  XNOR2_X1 U621 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U622 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n531) );
  INV_X1 U623 ( .A(G475), .ZN(n530) );
  INV_X1 U624 ( .A(n569), .ZN(n567) );
  NOR2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n618) );
  XNOR2_X1 U626 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n534) );
  XNOR2_X1 U627 ( .A(n535), .B(n534), .ZN(n773) );
  INV_X1 U628 ( .A(n773), .ZN(n549) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n716) );
  NOR2_X1 U630 ( .A1(n716), .A2(n728), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n536), .B(KEYINPUT108), .ZN(n538) );
  INV_X1 U632 ( .A(n560), .ZN(n537) );
  NAND2_X1 U633 ( .A1(n538), .A2(n537), .ZN(n541) );
  XNOR2_X1 U634 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n540) );
  INV_X1 U635 ( .A(KEYINPUT67), .ZN(n539) );
  AND2_X1 U636 ( .A1(n597), .A2(n729), .ZN(n542) );
  AND2_X1 U637 ( .A1(n374), .A2(n542), .ZN(n543) );
  XNOR2_X1 U638 ( .A(n543), .B(KEYINPUT81), .ZN(n544) );
  INV_X1 U639 ( .A(n729), .ZN(n613) );
  OR2_X1 U640 ( .A1(n731), .A2(n613), .ZN(n546) );
  NAND2_X1 U641 ( .A1(n549), .A2(n548), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n574), .A2(KEYINPUT44), .ZN(n572) );
  INV_X1 U643 ( .A(n597), .ZN(n550) );
  NOR2_X1 U644 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U645 ( .A1(n374), .A2(n729), .ZN(n553) );
  INV_X1 U646 ( .A(n554), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n555), .A2(n731), .ZN(n736) );
  NOR2_X1 U648 ( .A1(n736), .A2(n556), .ZN(n557) );
  XNOR2_X1 U649 ( .A(n557), .B(KEYINPUT31), .ZN(n706) );
  NAND2_X1 U650 ( .A1(n559), .A2(n726), .ZN(n580) );
  OR2_X1 U651 ( .A1(n560), .A2(n580), .ZN(n562) );
  INV_X1 U652 ( .A(KEYINPUT98), .ZN(n561) );
  XNOR2_X1 U653 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n563), .A2(n591), .ZN(n565) );
  INV_X1 U655 ( .A(KEYINPUT99), .ZN(n564) );
  INV_X1 U656 ( .A(n568), .ZN(n566) );
  NAND2_X1 U657 ( .A1(n567), .A2(n566), .ZN(n707) );
  NAND2_X1 U658 ( .A1(n707), .A2(n596), .ZN(n611) );
  XNOR2_X1 U659 ( .A(n570), .B(KEYINPUT109), .ZN(n571) );
  NAND2_X1 U660 ( .A1(n575), .A2(n358), .ZN(n577) );
  XNOR2_X1 U661 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n576) );
  NAND2_X1 U662 ( .A1(G953), .A2(G900), .ZN(n578) );
  NAND2_X1 U663 ( .A1(n579), .A2(n578), .ZN(n590) );
  OR2_X1 U664 ( .A1(n580), .A2(n588), .ZN(n581) );
  NOR2_X1 U665 ( .A1(n590), .A2(n581), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n731), .A2(n713), .ZN(n582) );
  XNOR2_X1 U667 ( .A(KEYINPUT30), .B(n582), .ZN(n620) );
  INV_X1 U668 ( .A(n620), .ZN(n583) );
  NOR2_X1 U669 ( .A1(n596), .A2(n626), .ZN(n587) );
  XNOR2_X1 U670 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n586) );
  XNOR2_X1 U671 ( .A(n587), .B(n586), .ZN(n772) );
  INV_X1 U672 ( .A(n588), .ZN(n714) );
  NOR2_X1 U673 ( .A1(n719), .A2(n716), .ZN(n589) );
  INV_X1 U674 ( .A(n749), .ZN(n739) );
  NOR2_X1 U675 ( .A1(n728), .A2(n590), .ZN(n614) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n614), .ZN(n594) );
  NAND2_X1 U677 ( .A1(n739), .A2(n605), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n592), .B(KEYINPUT42), .ZN(n593) );
  XNOR2_X1 U679 ( .A(KEYINPUT113), .B(n593), .ZN(n775) );
  INV_X1 U680 ( .A(n374), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n594), .A2(n613), .ZN(n599) );
  INV_X1 U682 ( .A(KEYINPUT110), .ZN(n595) );
  XNOR2_X1 U683 ( .A(n596), .B(n595), .ZN(n700) );
  INV_X1 U684 ( .A(n700), .ZN(n703) );
  NOR2_X1 U685 ( .A1(n597), .A2(n703), .ZN(n598) );
  NAND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n627) );
  XNOR2_X1 U687 ( .A(n701), .B(n608), .ZN(n610) );
  OR2_X1 U688 ( .A1(KEYINPUT47), .A2(n611), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n624) );
  INV_X1 U690 ( .A(n611), .ZN(n718) );
  NAND2_X1 U691 ( .A1(KEYINPUT47), .A2(n718), .ZN(n612) );
  XNOR2_X1 U692 ( .A(KEYINPUT85), .B(n612), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n631), .A2(n615), .ZN(n616) );
  AND2_X1 U695 ( .A1(n559), .A2(n616), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n699) );
  NOR2_X1 U698 ( .A1(n621), .A2(n699), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT83), .B(n622), .Z(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U701 ( .A1(n626), .A2(n707), .ZN(n711) );
  INV_X1 U702 ( .A(n711), .ZN(n633) );
  XOR2_X1 U703 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n630) );
  NOR2_X1 U704 ( .A1(n374), .A2(n627), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n628), .A2(n713), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n662) );
  NOR2_X1 U708 ( .A1(n638), .A2(KEYINPUT2), .ZN(n635) );
  OR2_X1 U709 ( .A1(n638), .A2(KEYINPUT88), .ZN(n636) );
  AND2_X1 U710 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(KEYINPUT88), .ZN(n639) );
  INV_X1 U712 ( .A(KEYINPUT66), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n679), .A2(G475), .ZN(n645) );
  XNOR2_X1 U714 ( .A(KEYINPUT92), .B(KEYINPUT124), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT59), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n647) );
  INV_X1 U718 ( .A(G952), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n646), .A2(G953), .ZN(n682) );
  NAND2_X1 U720 ( .A1(n679), .A2(G210), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U724 ( .A(G110), .B(KEYINPUT116), .Z(n653) );
  XNOR2_X1 U725 ( .A(n360), .B(n653), .ZN(G12) );
  XNOR2_X1 U726 ( .A(n654), .B(G119), .ZN(G21) );
  XNOR2_X1 U727 ( .A(n655), .B(G101), .ZN(G3) );
  NOR2_X1 U728 ( .A1(n660), .A2(n707), .ZN(n659) );
  XOR2_X1 U729 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n657) );
  XNOR2_X1 U730 ( .A(G107), .B(KEYINPUT26), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(G9) );
  NOR2_X1 U733 ( .A1(n660), .A2(n703), .ZN(n661) );
  XOR2_X1 U734 ( .A(G104), .B(n661), .Z(G6) );
  XNOR2_X1 U735 ( .A(n662), .B(G140), .ZN(G42) );
  NAND2_X1 U736 ( .A1(n679), .A2(G472), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT91), .B(KEYINPUT62), .Z(n663) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(n682), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(G57) );
  XOR2_X1 U743 ( .A(n671), .B(n670), .Z(n674) );
  XOR2_X1 U744 ( .A(n674), .B(n672), .Z(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(n762), .ZN(n678) );
  XNOR2_X1 U746 ( .A(G227), .B(n674), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n675), .A2(G900), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n676), .A2(G953), .ZN(n677) );
  NAND2_X1 U749 ( .A1(n678), .A2(n677), .ZN(G72) );
  NAND2_X1 U750 ( .A1(n687), .A2(G217), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(n683) );
  INV_X1 U752 ( .A(n682), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n683), .A2(n692), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n687), .A2(G478), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n686), .A2(n692), .ZN(G63) );
  NAND2_X1 U757 ( .A1(n687), .A2(G469), .ZN(n691) );
  XOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XOR2_X1 U759 ( .A(n689), .B(n688), .Z(n690) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(G54) );
  XOR2_X1 U762 ( .A(G128), .B(KEYINPUT117), .Z(n696) );
  INV_X1 U763 ( .A(n707), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n694), .A2(n701), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n696), .B(n695), .ZN(n698) );
  XOR2_X1 U766 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n697) );
  XNOR2_X1 U767 ( .A(n698), .B(n697), .ZN(G30) );
  XOR2_X1 U768 ( .A(G143), .B(n699), .Z(G45) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(G146), .ZN(G48) );
  NOR2_X1 U771 ( .A1(n703), .A2(n706), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G113), .B(KEYINPUT119), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n705), .B(n704), .ZN(G15) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U775 ( .A(G116), .B(n708), .Z(G18) );
  XNOR2_X1 U776 ( .A(G125), .B(n709), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(n711), .Z(G36) );
  NAND2_X1 U779 ( .A1(G952), .A2(n712), .ZN(n744) );
  NOR2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U782 ( .A(n717), .B(KEYINPUT120), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U785 ( .A(KEYINPUT121), .B(n722), .Z(n723) );
  NOR2_X1 U786 ( .A1(n750), .A2(n723), .ZN(n724) );
  XOR2_X1 U787 ( .A(KEYINPUT122), .B(n724), .Z(n741) );
  NOR2_X1 U788 ( .A1(n726), .A2(n374), .ZN(n727) );
  XOR2_X1 U789 ( .A(KEYINPUT50), .B(n727), .Z(n734) );
  NAND2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U791 ( .A(n730), .B(KEYINPUT49), .ZN(n732) );
  NOR2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U795 ( .A(KEYINPUT51), .B(n737), .Z(n738) );
  NAND2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U798 ( .A(KEYINPUT52), .B(n742), .Z(n743) );
  NOR2_X1 U799 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U800 ( .A(KEYINPUT123), .B(n745), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n746), .A2(KEYINPUT84), .ZN(n747) );
  XNOR2_X1 U802 ( .A(n747), .B(KEYINPUT87), .ZN(n748) );
  XNOR2_X1 U803 ( .A(n748), .B(KEYINPUT2), .ZN(n752) );
  NOR2_X1 U804 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n756), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U808 ( .A(n757), .B(G101), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n761) );
  NOR2_X1 U810 ( .A1(n762), .A2(G898), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n771) );
  AND2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n769) );
  INV_X1 U813 ( .A(G898), .ZN(n767) );
  NAND2_X1 U814 ( .A1(G224), .A2(G953), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n764), .B(KEYINPUT61), .ZN(n765) );
  XNOR2_X1 U816 ( .A(n765), .B(KEYINPUT125), .ZN(n766) );
  NOR2_X1 U817 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U818 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U819 ( .A(n771), .B(n770), .Z(G69) );
  XOR2_X1 U820 ( .A(G131), .B(n772), .Z(G33) );
  XOR2_X1 U821 ( .A(G122), .B(KEYINPUT126), .Z(n774) );
  XNOR2_X1 U822 ( .A(n773), .B(n774), .ZN(G24) );
  XOR2_X1 U823 ( .A(n775), .B(G137), .Z(G39) );
endmodule

