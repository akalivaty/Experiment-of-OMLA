

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731;

  AND2_X1 U369 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U370 ( .A(n487), .B(n486), .ZN(n514) );
  NAND2_X1 U371 ( .A1(n537), .A2(n484), .ZN(n487) );
  XNOR2_X1 U372 ( .A(n478), .B(n477), .ZN(n528) );
  NAND2_X1 U373 ( .A1(n349), .A2(n348), .ZN(n562) );
  XNOR2_X1 U374 ( .A(n464), .B(n350), .ZN(n349) );
  INV_X1 U375 ( .A(n468), .ZN(n348) );
  OR2_X1 U376 ( .A1(n592), .A2(n590), .ZN(n464) );
  INV_X1 U377 ( .A(n463), .ZN(n350) );
  XNOR2_X1 U378 ( .A(n368), .B(G101), .ZN(n398) );
  INV_X1 U379 ( .A(G953), .ZN(n724) );
  NOR2_X2 U380 ( .A1(n619), .A2(n603), .ZN(n607) );
  AND2_X2 U381 ( .A1(n514), .A2(n631), .ZN(n534) );
  NAND2_X1 U382 ( .A1(n528), .A2(n479), .ZN(n481) );
  XNOR2_X1 U383 ( .A(KEYINPUT3), .B(G119), .ZN(n402) );
  NAND2_X1 U384 ( .A1(n566), .A2(n664), .ZN(n642) );
  XNOR2_X2 U385 ( .A(n558), .B(KEYINPUT112), .ZN(n637) );
  NOR2_X2 U386 ( .A1(n681), .A2(n523), .ZN(n504) );
  XNOR2_X1 U387 ( .A(n562), .B(KEYINPUT19), .ZN(n351) );
  XNOR2_X1 U388 ( .A(n464), .B(n463), .ZN(n352) );
  XNOR2_X1 U389 ( .A(n562), .B(KEYINPUT19), .ZN(n576) );
  BUF_X1 U390 ( .A(n619), .Z(n690) );
  XNOR2_X2 U391 ( .A(n381), .B(G140), .ZN(n714) );
  XNOR2_X2 U392 ( .A(n716), .B(G146), .ZN(n407) );
  XNOR2_X2 U393 ( .A(n421), .B(n367), .ZN(n716) );
  INV_X1 U394 ( .A(n728), .ZN(n539) );
  INV_X1 U395 ( .A(KEYINPUT102), .ZN(n432) );
  XNOR2_X1 U396 ( .A(n548), .B(n547), .ZN(n652) );
  XNOR2_X1 U397 ( .A(n442), .B(G475), .ZN(n443) );
  XNOR2_X1 U398 ( .A(n552), .B(n483), .ZN(n500) );
  XNOR2_X1 U399 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U400 ( .A(n370), .B(n369), .ZN(n371) );
  NOR2_X1 U401 ( .A1(n527), .A2(n417), .ZN(n555) );
  OR2_X1 U402 ( .A1(n697), .A2(G902), .ZN(n395) );
  XNOR2_X1 U403 ( .A(n598), .B(n597), .ZN(n699) );
  XOR2_X1 U404 ( .A(n384), .B(KEYINPUT23), .Z(n353) );
  AND2_X1 U405 ( .A1(n583), .A2(n582), .ZN(n354) );
  OR2_X1 U406 ( .A1(n580), .A2(n579), .ZN(n355) );
  NOR2_X1 U407 ( .A1(n533), .A2(n532), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n448), .B(n371), .ZN(n373) );
  XNOR2_X1 U409 ( .A(KEYINPUT28), .B(n551), .ZN(n357) );
  XOR2_X1 U410 ( .A(KEYINPUT30), .B(n411), .Z(n358) );
  XOR2_X1 U411 ( .A(n394), .B(n393), .Z(n359) );
  XNOR2_X1 U412 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n444), .B(n443), .ZN(n489) );
  NOR2_X1 U414 ( .A1(n581), .A2(n355), .ZN(n582) );
  XNOR2_X1 U415 ( .A(G137), .B(G110), .ZN(n384) );
  XNOR2_X1 U416 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U417 ( .A(n434), .B(n714), .ZN(n441) );
  INV_X1 U418 ( .A(KEYINPUT114), .ZN(n547) );
  INV_X1 U419 ( .A(G469), .ZN(n375) );
  NOR2_X1 U420 ( .A1(n588), .A2(n587), .ZN(n721) );
  XNOR2_X1 U421 ( .A(n385), .B(n353), .ZN(n386) );
  XNOR2_X1 U422 ( .A(KEYINPUT36), .B(KEYINPUT88), .ZN(n564) );
  BUF_X1 U423 ( .A(n721), .Z(n722) );
  XNOR2_X1 U424 ( .A(n565), .B(n564), .ZN(n566) );
  INV_X2 U425 ( .A(G143), .ZN(n466) );
  XNOR2_X2 U426 ( .A(n466), .B(G128), .ZN(n452) );
  INV_X1 U427 ( .A(n452), .ZN(n361) );
  NAND2_X1 U428 ( .A1(G134), .A2(n361), .ZN(n364) );
  INV_X1 U429 ( .A(G134), .ZN(n362) );
  NAND2_X1 U430 ( .A1(n362), .A2(n452), .ZN(n363) );
  NAND2_X1 U431 ( .A1(n364), .A2(n363), .ZN(n421) );
  XOR2_X1 U432 ( .A(KEYINPUT4), .B(G131), .Z(n366) );
  XNOR2_X1 U433 ( .A(KEYINPUT72), .B(G137), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n367) );
  INV_X1 U435 ( .A(KEYINPUT70), .ZN(n368) );
  XNOR2_X1 U436 ( .A(G110), .B(G104), .ZN(n700) );
  XNOR2_X1 U437 ( .A(n398), .B(n700), .ZN(n448) );
  NAND2_X1 U438 ( .A1(G227), .A2(n724), .ZN(n370) );
  INV_X1 U439 ( .A(KEYINPUT97), .ZN(n369) );
  XOR2_X1 U440 ( .A(G107), .B(G140), .Z(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n407), .B(n374), .ZN(n621) );
  NOR2_X2 U443 ( .A1(G902), .A2(n621), .ZN(n376) );
  XNOR2_X2 U444 ( .A(n376), .B(n375), .ZN(n552) );
  XNOR2_X1 U445 ( .A(KEYINPUT15), .B(G902), .ZN(n460) );
  NAND2_X1 U446 ( .A1(G234), .A2(n460), .ZN(n377) );
  XNOR2_X1 U447 ( .A(KEYINPUT20), .B(n377), .ZN(n391) );
  AND2_X1 U448 ( .A1(n391), .A2(G221), .ZN(n379) );
  INV_X1 U449 ( .A(KEYINPUT21), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n659) );
  INV_X1 U451 ( .A(G146), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n380), .B(G125), .ZN(n446) );
  XNOR2_X1 U453 ( .A(n446), .B(KEYINPUT10), .ZN(n381) );
  XOR2_X1 U454 ( .A(G128), .B(G119), .Z(n383) );
  XOR2_X1 U455 ( .A(KEYINPUT24), .B(KEYINPUT98), .Z(n382) );
  XNOR2_X1 U456 ( .A(n714), .B(n386), .ZN(n390) );
  NAND2_X1 U457 ( .A1(n724), .A2(G234), .ZN(n388) );
  XNOR2_X1 U458 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n422) );
  NAND2_X1 U460 ( .A1(G221), .A2(n422), .ZN(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n697) );
  NAND2_X1 U462 ( .A1(n391), .A2(G217), .ZN(n394) );
  XNOR2_X1 U463 ( .A(KEYINPUT25), .B(KEYINPUT79), .ZN(n392) );
  XNOR2_X1 U464 ( .A(n392), .B(KEYINPUT78), .ZN(n393) );
  XNOR2_X2 U465 ( .A(n395), .B(n359), .ZN(n658) );
  NOR2_X2 U466 ( .A1(n659), .A2(n658), .ZN(n665) );
  NAND2_X1 U467 ( .A1(n552), .A2(n665), .ZN(n527) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n396) );
  XOR2_X1 U469 ( .A(KEYINPUT77), .B(n396), .Z(n435) );
  NAND2_X1 U470 ( .A1(n435), .A2(G210), .ZN(n400) );
  XNOR2_X1 U471 ( .A(G116), .B(KEYINPUT99), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n405) );
  INV_X1 U474 ( .A(G113), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n455) );
  XOR2_X1 U476 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n403) );
  XNOR2_X1 U477 ( .A(n455), .B(n403), .ZN(n404) );
  XNOR2_X1 U478 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n407), .B(n406), .ZN(n605) );
  INV_X1 U480 ( .A(G902), .ZN(n427) );
  NAND2_X1 U481 ( .A1(n605), .A2(n427), .ZN(n408) );
  INV_X1 U482 ( .A(G472), .ZN(n603) );
  XNOR2_X2 U483 ( .A(n408), .B(n603), .ZN(n661) );
  INV_X1 U484 ( .A(n661), .ZN(n526) );
  NOR2_X1 U485 ( .A1(G237), .A2(G902), .ZN(n409) );
  XNOR2_X1 U486 ( .A(n409), .B(KEYINPUT76), .ZN(n461) );
  INV_X1 U487 ( .A(G214), .ZN(n410) );
  OR2_X1 U488 ( .A1(n461), .A2(n410), .ZN(n646) );
  NAND2_X1 U489 ( .A1(n526), .A2(n646), .ZN(n411) );
  NAND2_X1 U490 ( .A1(G234), .A2(G237), .ZN(n412) );
  XNOR2_X1 U491 ( .A(n412), .B(KEYINPUT14), .ZN(n414) );
  NAND2_X1 U492 ( .A1(G902), .A2(n414), .ZN(n469) );
  NOR2_X1 U493 ( .A1(G900), .A2(n469), .ZN(n413) );
  NAND2_X1 U494 ( .A1(G953), .A2(n413), .ZN(n416) );
  NAND2_X1 U495 ( .A1(G952), .A2(n414), .ZN(n415) );
  XNOR2_X1 U496 ( .A(KEYINPUT95), .B(n415), .ZN(n677) );
  NAND2_X1 U497 ( .A1(n677), .A2(n724), .ZN(n473) );
  NAND2_X1 U498 ( .A1(n416), .A2(n473), .ZN(n492) );
  NAND2_X1 U499 ( .A1(n358), .A2(n492), .ZN(n417) );
  XOR2_X1 U500 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n419) );
  XNOR2_X1 U501 ( .A(KEYINPUT108), .B(KEYINPUT9), .ZN(n418) );
  XNOR2_X1 U502 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U503 ( .A(n421), .B(n420), .Z(n424) );
  NAND2_X1 U504 ( .A1(G217), .A2(n422), .ZN(n423) );
  XNOR2_X1 U505 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U506 ( .A(G122), .B(G116), .ZN(n425) );
  XNOR2_X1 U507 ( .A(n425), .B(G107), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n426), .B(n457), .ZN(n691) );
  NAND2_X1 U509 ( .A1(n691), .A2(n427), .ZN(n428) );
  INV_X1 U510 ( .A(G478), .ZN(n689) );
  XNOR2_X1 U511 ( .A(n428), .B(n689), .ZN(n490) );
  XOR2_X1 U512 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n430) );
  XNOR2_X1 U513 ( .A(G113), .B(KEYINPUT103), .ZN(n429) );
  XNOR2_X1 U514 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U515 ( .A(n431), .B(KEYINPUT104), .ZN(n433) );
  XNOR2_X1 U516 ( .A(G143), .B(G131), .ZN(n439) );
  NAND2_X1 U517 ( .A1(G214), .A2(n435), .ZN(n437) );
  XOR2_X1 U518 ( .A(G104), .B(G122), .Z(n436) );
  XNOR2_X1 U519 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U520 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U521 ( .A(n441), .B(n440), .ZN(n612) );
  NOR2_X1 U522 ( .A1(n612), .A2(G902), .ZN(n444) );
  XNOR2_X1 U523 ( .A(KEYINPUT105), .B(KEYINPUT13), .ZN(n442) );
  NOR2_X1 U524 ( .A1(n490), .A2(n489), .ZN(n505) );
  NAND2_X1 U525 ( .A1(n555), .A2(n505), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n445) );
  XNOR2_X1 U527 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U528 ( .A(n448), .B(n447), .ZN(n454) );
  XNOR2_X1 U529 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n450) );
  NAND2_X1 U530 ( .A1(n724), .A2(G224), .ZN(n449) );
  XNOR2_X1 U531 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U532 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U533 ( .A(n454), .B(n453), .ZN(n459) );
  INV_X1 U534 ( .A(n455), .ZN(n456) );
  XNOR2_X1 U535 ( .A(n456), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U536 ( .A(n458), .B(n457), .ZN(n702) );
  XNOR2_X1 U537 ( .A(n459), .B(n702), .ZN(n592) );
  INV_X1 U538 ( .A(n460), .ZN(n590) );
  INV_X1 U539 ( .A(G210), .ZN(n591) );
  OR2_X1 U540 ( .A1(n461), .A2(n591), .ZN(n462) );
  XNOR2_X1 U541 ( .A(n462), .B(KEYINPUT94), .ZN(n463) );
  NOR2_X1 U542 ( .A1(n465), .A2(n352), .ZN(n579) );
  XNOR2_X1 U543 ( .A(n579), .B(n466), .ZN(G45) );
  AND2_X1 U544 ( .A1(n489), .A2(n490), .ZN(n645) );
  INV_X1 U545 ( .A(n659), .ZN(n467) );
  AND2_X1 U546 ( .A1(n645), .A2(n467), .ZN(n479) );
  INV_X1 U547 ( .A(n646), .ZN(n468) );
  INV_X1 U548 ( .A(n469), .ZN(n470) );
  NOR2_X1 U549 ( .A1(G898), .A2(n724), .ZN(n703) );
  NAND2_X1 U550 ( .A1(n470), .A2(n703), .ZN(n471) );
  XNOR2_X1 U551 ( .A(n471), .B(KEYINPUT96), .ZN(n472) );
  NAND2_X1 U552 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U553 ( .A1(n576), .A2(n474), .ZN(n478) );
  XNOR2_X1 U554 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n476) );
  INV_X1 U555 ( .A(KEYINPUT69), .ZN(n475) );
  XNOR2_X1 U556 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U557 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n480) );
  XNOR2_X1 U558 ( .A(n481), .B(n480), .ZN(n513) );
  XNOR2_X1 U559 ( .A(KEYINPUT110), .B(KEYINPUT6), .ZN(n482) );
  XNOR2_X1 U560 ( .A(n661), .B(n482), .ZN(n502) );
  NOR2_X2 U561 ( .A1(n513), .A2(n502), .ZN(n537) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(KEYINPUT67), .Z(n483) );
  INV_X1 U563 ( .A(n500), .ZN(n511) );
  INV_X1 U564 ( .A(n658), .ZN(n491) );
  NOR2_X1 U565 ( .A1(n511), .A2(n491), .ZN(n484) );
  XNOR2_X1 U566 ( .A(KEYINPUT81), .B(KEYINPUT32), .ZN(n485) );
  XNOR2_X1 U567 ( .A(n485), .B(KEYINPUT65), .ZN(n486) );
  XOR2_X1 U568 ( .A(G119), .B(KEYINPUT127), .Z(n488) );
  XNOR2_X1 U569 ( .A(n514), .B(n488), .ZN(G21) );
  INV_X1 U570 ( .A(n511), .ZN(n664) );
  XNOR2_X1 U571 ( .A(KEYINPUT106), .B(n489), .ZN(n519) );
  INV_X1 U572 ( .A(n490), .ZN(n518) );
  NOR2_X2 U573 ( .A1(n519), .A2(n518), .ZN(n558) );
  NOR2_X1 U574 ( .A1(n491), .A2(n659), .ZN(n493) );
  NAND2_X1 U575 ( .A1(n493), .A2(n492), .ZN(n550) );
  INV_X1 U576 ( .A(n550), .ZN(n494) );
  AND2_X1 U577 ( .A1(n502), .A2(n494), .ZN(n495) );
  AND2_X1 U578 ( .A1(n637), .A2(n495), .ZN(n561) );
  NAND2_X1 U579 ( .A1(n561), .A2(n646), .ZN(n496) );
  NOR2_X1 U580 ( .A1(n664), .A2(n496), .ZN(n498) );
  XNOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n497) );
  XNOR2_X1 U582 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U583 ( .A1(n499), .A2(n352), .ZN(n586) );
  XNOR2_X1 U584 ( .A(n586), .B(G140), .ZN(G42) );
  NAND2_X1 U585 ( .A1(n500), .A2(n665), .ZN(n501) );
  XNOR2_X1 U586 ( .A(n501), .B(KEYINPUT75), .ZN(n521) );
  AND2_X2 U587 ( .A1(n521), .A2(n502), .ZN(n503) );
  XNOR2_X2 U588 ( .A(n503), .B(KEYINPUT33), .ZN(n681) );
  INV_X1 U589 ( .A(n528), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n504), .B(KEYINPUT34), .ZN(n507) );
  XNOR2_X1 U591 ( .A(n505), .B(KEYINPUT80), .ZN(n506) );
  NAND2_X1 U592 ( .A1(n507), .A2(n506), .ZN(n509) );
  XNOR2_X1 U593 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U594 ( .A(n509), .B(n508), .ZN(n729) );
  NOR2_X1 U595 ( .A1(n729), .A2(KEYINPUT44), .ZN(n515) );
  AND2_X1 U596 ( .A1(n658), .A2(n661), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n511), .A2(n510), .ZN(n512) );
  OR2_X1 U598 ( .A1(n513), .A2(n512), .ZN(n631) );
  NAND2_X1 U599 ( .A1(n515), .A2(n534), .ZN(n516) );
  XNOR2_X1 U600 ( .A(KEYINPUT74), .B(n516), .ZN(n517) );
  INV_X1 U601 ( .A(n517), .ZN(n543) );
  AND2_X1 U602 ( .A1(n729), .A2(KEYINPUT44), .ZN(n533) );
  NAND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U604 ( .A(n520), .B(KEYINPUT109), .ZN(n639) );
  NOR2_X1 U605 ( .A1(n558), .A2(n639), .ZN(n574) );
  XNOR2_X1 U606 ( .A(n574), .B(KEYINPUT82), .ZN(n531) );
  BUF_X1 U607 ( .A(n521), .Z(n522) );
  NAND2_X1 U608 ( .A1(n522), .A2(n526), .ZN(n670) );
  NOR2_X1 U609 ( .A1(n670), .A2(n523), .ZN(n525) );
  XNOR2_X1 U610 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n524) );
  XNOR2_X1 U611 ( .A(n525), .B(n524), .ZN(n640) );
  NOR2_X1 U612 ( .A1(n527), .A2(n526), .ZN(n529) );
  AND2_X1 U613 ( .A1(n529), .A2(n528), .ZN(n626) );
  NOR2_X1 U614 ( .A1(n640), .A2(n626), .ZN(n530) );
  NOR2_X1 U615 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U616 ( .A(n534), .ZN(n535) );
  NAND2_X1 U617 ( .A1(n535), .A2(KEYINPUT44), .ZN(n540) );
  NOR2_X1 U618 ( .A1(n664), .A2(n658), .ZN(n536) );
  NAND2_X1 U619 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U620 ( .A(n538), .B(KEYINPUT111), .ZN(n728) );
  NAND2_X1 U621 ( .A1(n356), .A2(n541), .ZN(n542) );
  NOR2_X2 U622 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U623 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n544) );
  XNOR2_X1 U624 ( .A(n545), .B(n544), .ZN(n705) );
  XNOR2_X1 U625 ( .A(n352), .B(KEYINPUT38), .ZN(n647) );
  NAND2_X1 U626 ( .A1(n647), .A2(n646), .ZN(n548) );
  NAND2_X1 U627 ( .A1(n652), .A2(n645), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n549), .B(KEYINPUT41), .ZN(n680) );
  NOR2_X1 U629 ( .A1(n661), .A2(n550), .ZN(n551) );
  NAND2_X1 U630 ( .A1(n357), .A2(n552), .ZN(n575) );
  INV_X1 U631 ( .A(n575), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n680), .A2(n553), .ZN(n554) );
  XNOR2_X1 U633 ( .A(KEYINPUT42), .B(n554), .ZN(n730) );
  XOR2_X1 U634 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n557) );
  NAND2_X1 U635 ( .A1(n555), .A2(n647), .ZN(n556) );
  XNOR2_X1 U636 ( .A(n557), .B(n556), .ZN(n585) );
  NAND2_X1 U637 ( .A1(n558), .A2(n585), .ZN(n559) );
  XNOR2_X1 U638 ( .A(KEYINPUT40), .B(n559), .ZN(n731) );
  AND2_X1 U639 ( .A1(n730), .A2(n731), .ZN(n560) );
  XNOR2_X1 U640 ( .A(n560), .B(n360), .ZN(n583) );
  XNOR2_X1 U641 ( .A(n561), .B(KEYINPUT115), .ZN(n563) );
  NOR2_X1 U642 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U643 ( .A(n642), .B(KEYINPUT86), .ZN(n573) );
  INV_X1 U644 ( .A(KEYINPUT47), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n553), .A2(n351), .ZN(n632) );
  NOR2_X1 U646 ( .A1(n574), .A2(n632), .ZN(n569) );
  NAND2_X1 U647 ( .A1(n569), .A2(KEYINPUT82), .ZN(n567) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n569), .A2(KEYINPUT47), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n573), .A2(n572), .ZN(n581) );
  INV_X1 U652 ( .A(n574), .ZN(n651) );
  NOR2_X1 U653 ( .A1(n575), .A2(KEYINPUT82), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n577), .A2(n351), .ZN(n578) );
  NOR2_X1 U655 ( .A1(n651), .A2(n578), .ZN(n580) );
  XNOR2_X1 U656 ( .A(KEYINPUT48), .B(KEYINPUT73), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n354), .B(n584), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n585), .A2(n639), .ZN(n644) );
  NAND2_X1 U659 ( .A1(n586), .A2(n644), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n705), .A2(n721), .ZN(n589) );
  XNOR2_X2 U661 ( .A(n589), .B(KEYINPUT2), .ZN(n679) );
  NAND2_X2 U662 ( .A1(n679), .A2(n590), .ZN(n619) );
  NOR2_X1 U663 ( .A1(n619), .A2(n591), .ZN(n595) );
  XNOR2_X1 U664 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n593) );
  XNOR2_X1 U665 ( .A(n592), .B(n593), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n595), .B(n594), .ZN(n599) );
  INV_X1 U667 ( .A(G952), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n596), .A2(G953), .ZN(n598) );
  INV_X1 U669 ( .A(KEYINPUT92), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n599), .A2(n699), .ZN(n602) );
  XNOR2_X1 U671 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT85), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n602), .B(n601), .ZN(G51) );
  INV_X1 U674 ( .A(KEYINPUT63), .ZN(n610) );
  XNOR2_X1 U675 ( .A(KEYINPUT90), .B(KEYINPUT62), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n608), .A2(n699), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(G57) );
  INV_X1 U680 ( .A(n619), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n611), .A2(G475), .ZN(n615) );
  XNOR2_X1 U682 ( .A(KEYINPUT91), .B(KEYINPUT59), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n612), .B(n613), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X2 U685 ( .A1(n616), .A2(n699), .ZN(n618) );
  XNOR2_X1 U686 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(G60) );
  INV_X1 U688 ( .A(n690), .ZN(n695) );
  NAND2_X1 U689 ( .A1(n695), .A2(G469), .ZN(n623) );
  XOR2_X1 U690 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U693 ( .A1(n624), .A2(n699), .ZN(G54) );
  NAND2_X1 U694 ( .A1(n637), .A2(n626), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(G104), .ZN(G6) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT27), .ZN(n630) );
  XOR2_X1 U697 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U698 ( .A1(n626), .A2(n639), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G9) );
  XNOR2_X1 U701 ( .A(G110), .B(n631), .ZN(G12) );
  XOR2_X1 U702 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  INV_X1 U703 ( .A(n632), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n639), .A2(n635), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G30) );
  NAND2_X1 U706 ( .A1(n637), .A2(n635), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n637), .A2(n640), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(G113), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(G116), .ZN(G18) );
  XOR2_X1 U712 ( .A(G125), .B(KEYINPUT37), .Z(n643) );
  XNOR2_X1 U713 ( .A(n642), .B(n643), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n644), .ZN(G36) );
  INV_X1 U715 ( .A(n681), .ZN(n657) );
  INV_X1 U716 ( .A(n645), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U719 ( .A(KEYINPUT118), .B(n650), .Z(n654) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U722 ( .A(KEYINPUT119), .B(n655), .Z(n656) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n674) );
  NAND2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n660), .Z(n662) );
  NAND2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U727 ( .A(KEYINPUT117), .B(n663), .ZN(n668) );
  NOR2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U729 ( .A(KEYINPUT50), .B(n666), .Z(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  NAND2_X1 U733 ( .A1(n680), .A2(n672), .ZN(n673) );
  NAND2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n675), .B(KEYINPUT120), .ZN(n676) );
  XNOR2_X1 U736 ( .A(KEYINPUT52), .B(n676), .ZN(n678) );
  NAND2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n687) );
  BUF_X1 U738 ( .A(n679), .Z(n685) );
  INV_X1 U739 ( .A(n680), .ZN(n682) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  OR2_X1 U741 ( .A1(n683), .A2(G953), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U744 ( .A(KEYINPUT53), .B(n688), .Z(G75) );
  NOR2_X1 U745 ( .A1(n690), .A2(n689), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n691), .B(KEYINPUT122), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U748 ( .A1(n699), .A2(n694), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n695), .A2(G217), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n699), .A2(n698), .ZN(G66) );
  XNOR2_X1 U752 ( .A(n700), .B(G101), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n712) );
  NAND2_X1 U755 ( .A1(n705), .A2(n724), .ZN(n710) );
  XOR2_X1 U756 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n707) );
  NAND2_X1 U757 ( .A1(G224), .A2(G953), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U759 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U762 ( .A(KEYINPUT124), .B(n713), .ZN(G69) );
  XOR2_X1 U763 ( .A(n714), .B(KEYINPUT97), .Z(n715) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n723) );
  XNOR2_X1 U765 ( .A(n723), .B(KEYINPUT125), .ZN(n717) );
  XNOR2_X1 U766 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(G900), .A2(n718), .ZN(n719) );
  NAND2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n720), .B(KEYINPUT126), .ZN(n727) );
  XNOR2_X1 U770 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n727), .A2(n726), .ZN(G72) );
  XOR2_X1 U773 ( .A(G101), .B(n728), .Z(G3) );
  XOR2_X1 U774 ( .A(n729), .B(G122), .Z(G24) );
  XNOR2_X1 U775 ( .A(G137), .B(n730), .ZN(G39) );
  XNOR2_X1 U776 ( .A(G131), .B(n731), .ZN(G33) );
endmodule

