//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n467), .B2(KEYINPUT67), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT67), .B(G125), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n475), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(new_n470), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n466), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n484), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n475), .A2(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n469), .B2(new_n470), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n496), .C1(new_n470), .C2(new_n469), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n474), .A2(new_n505), .A3(new_n496), .A4(new_n499), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n497), .A2(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  AND2_X1   g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n474), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n474), .B2(new_n509), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n475), .A2(G114), .ZN(new_n513));
  OAI21_X1  g088(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G164));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(G50), .A2(new_n525), .B1(new_n530), .B2(G88), .ZN(new_n531));
  INV_X1    g106(.A(G75), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  OR3_X1    g108(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT75), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT75), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(G62), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(KEYINPUT74), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n531), .A2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n525), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n547));
  AND2_X1   g122(.A1(G63), .A2(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n546), .A2(new_n547), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(new_n528), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n517), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  AOI22_X1  g133(.A1(G52), .A2(new_n525), .B1(new_n530), .B2(G90), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(new_n530), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n525), .A2(G43), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n517), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI211_X1 g149(.A(KEYINPUT78), .B(new_n573), .C1(new_n524), .C2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(KEYINPUT79), .B(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n528), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(G78), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n518), .A2(new_n521), .B1(KEYINPUT6), .B2(new_n517), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT78), .B(KEYINPUT9), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n581), .A2(G53), .A3(G543), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(G91), .A3(new_n528), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n575), .A2(new_n580), .A3(new_n583), .A4(new_n584), .ZN(G299));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n517), .B1(new_n553), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n522), .A2(new_n523), .ZN(new_n588));
  NAND2_X1  g163(.A1(G49), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT81), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n581), .A2(new_n591), .A3(G49), .A4(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n529), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n581), .A2(KEYINPUT80), .A3(G87), .A4(new_n528), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(KEYINPUT82), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT82), .B1(new_n593), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(G288));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n526), .B2(new_n527), .ZN(new_n603));
  AND2_X1   g178(.A1(G73), .A2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n522), .A2(G86), .A3(new_n528), .A4(new_n523), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n523), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n530), .A2(G85), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n525), .A2(G47), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n517), .C2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n553), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n525), .A2(G54), .B1(new_n615), .B2(G651), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n529), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n529), .B2(new_n617), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n616), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G171), .B2(new_n622), .ZN(G284));
  XOR2_X1   g199(.A(G284), .B(KEYINPUT84), .Z(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n622), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n622), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G168), .B2(new_n622), .ZN(G280));
  INV_X1    g203(.A(new_n621), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n566), .A2(new_n622), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n621), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n637), .B1(new_n488), .B2(new_n638), .C1(new_n639), .C2(new_n491), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n474), .A2(new_n477), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT85), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n642), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT87), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n659), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n668), .B(KEYINPUT17), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n666), .C1(new_n676), .C2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n670), .A3(new_n665), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n685), .A2(KEYINPUT20), .A3(new_n688), .ZN(new_n694));
  OAI221_X1 g269(.A(new_n690), .B1(new_n688), .B2(new_n689), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G168), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT97), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G1966), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(G1966), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n710), .B(new_n711), .C1(G2090), .C2(new_n715), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n715), .A2(KEYINPUT99), .A3(G2090), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n712), .A2(G32), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n721), .A2(new_n722), .B1(G105), .B2(new_n477), .ZN(new_n723));
  INV_X1    g298(.A(G141), .ZN(new_n724));
  INV_X1    g299(.A(G129), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n723), .B1(new_n488), .B2(new_n724), .C1(new_n725), .C2(new_n491), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n718), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT27), .ZN(new_n728));
  INV_X1    g303(.A(G1996), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT99), .B1(new_n715), .B2(G2090), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n717), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n706), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n706), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT98), .Z(new_n736));
  NAND2_X1  g311(.A1(G160), .A2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(new_n712), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT96), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(G299), .A2(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n706), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT23), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n736), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n629), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G4), .B2(G16), .ZN(new_n751));
  INV_X1    g326(.A(G1348), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n712), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  INV_X1    g333(.A(G128), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n757), .B1(new_n488), .B2(new_n758), .C1(new_n759), .C2(new_n491), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n751), .A2(new_n752), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n753), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n706), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n567), .B2(new_n706), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1341), .Z(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G1961), .B2(new_n734), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n712), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n712), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT30), .B(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n712), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n640), .B2(new_n712), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n712), .A2(G33), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G139), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n780), .B1(new_n475), .B2(new_n781), .C1(new_n488), .C2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(new_n712), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n777), .B1(new_n785), .B2(G2072), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n772), .B(new_n786), .C1(G2072), .C2(new_n785), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n764), .A2(new_n768), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n716), .A2(new_n732), .A3(new_n749), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n706), .A2(G23), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n593), .A2(new_n598), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n706), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n792), .B(new_n793), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT95), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n706), .A2(G22), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G303), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1971), .ZN(new_n802));
  MUX2_X1   g377(.A(G6), .B(G305), .S(G16), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NAND4_X1  g380(.A1(new_n797), .A2(new_n799), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n712), .A2(G25), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n812));
  INV_X1    g387(.A(G131), .ZN(new_n813));
  INV_X1    g388(.A(G119), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n488), .B2(new_n813), .C1(new_n814), .C2(new_n491), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT94), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT94), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  MUX2_X1   g397(.A(G24), .B(G290), .S(G16), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1986), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n807), .A2(new_n808), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n807), .A2(new_n828), .A3(new_n808), .A4(new_n825), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n789), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT100), .ZN(G311));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(G150));
  NAND2_X1  g408(.A1(new_n530), .A2(G93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n525), .A2(G55), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n834), .B(new_n835), .C1(new_n517), .C2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n566), .A3(new_n840), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n837), .A2(new_n566), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n621), .A2(new_n630), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n847), .A2(new_n848), .A3(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n837), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n640), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n726), .B(G164), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(new_n783), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n783), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n760), .B(KEYINPUT103), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(G142), .B(new_n475), .C1(new_n486), .C2(new_n487), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n475), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n861), .B1(new_n862), .B2(new_n491), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n644), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n818), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n857), .B2(new_n858), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n860), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n860), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n855), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n855), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(new_n870), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n853), .B(new_n871), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(G395));
  NAND2_X1  g453(.A1(new_n837), .A2(new_n622), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n791), .B(G290), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n593), .A2(new_n598), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G290), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT108), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(G305), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(KEYINPUT109), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n621), .B(G299), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n633), .B(KEYINPUT106), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n843), .Z(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n893), .B2(new_n900), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n892), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n879), .B1(new_n903), .B2(new_n622), .ZN(G295));
  OAI21_X1  g479(.A(new_n879), .B1(new_n903), .B2(new_n622), .ZN(G331));
  NAND2_X1  g480(.A1(G171), .A2(G168), .ZN(new_n906));
  NAND2_X1  g481(.A1(G301), .A2(G286), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n843), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n841), .A2(new_n906), .A3(new_n842), .A4(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n894), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(KEYINPUT110), .C1(new_n893), .C2(new_n911), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n891), .B(new_n913), .C1(KEYINPUT110), .C2(new_n912), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n889), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n911), .A2(new_n893), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n898), .B2(new_n911), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n914), .A2(KEYINPUT43), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT43), .B1(new_n921), .B2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT44), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n914), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n921), .B2(new_n919), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n927), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n507), .B2(new_n515), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n473), .A2(G40), .A3(new_n480), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n818), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(new_n820), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n760), .B(G2067), .Z(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n726), .B(G1996), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n820), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(G290), .B(G1986), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n933), .B1(new_n930), .B2(KEYINPUT50), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n946), .B(new_n929), .C1(new_n507), .C2(new_n515), .ZN(new_n947));
  AOI21_X1  g522(.A(G1961), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n513), .A2(new_n514), .ZN(new_n950));
  INV_X1    g525(.A(new_n512), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n510), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n495), .A2(KEYINPUT71), .A3(new_n496), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n501), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n504), .A2(new_n506), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT45), .B1(new_n957), .B2(new_n929), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n931), .A2(G1384), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n507), .B2(new_n515), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT67), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n485), .B2(new_n464), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n471), .A3(new_n463), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n961), .B(new_n479), .C1(new_n964), .C2(G2105), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(KEYINPUT53), .A3(new_n771), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT111), .B1(new_n958), .B2(new_n966), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n933), .B1(new_n957), .B2(new_n959), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n932), .ZN(new_n972));
  AOI21_X1  g547(.A(G2078), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n949), .B(new_n968), .C1(new_n973), .C2(KEYINPUT53), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT126), .B1(new_n974), .B2(G171), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n958), .A2(new_n966), .A3(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n971), .B1(new_n970), .B2(new_n932), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n771), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n948), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT126), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n981), .A3(G301), .A4(new_n968), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n949), .B1(new_n973), .B2(KEYINPUT53), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n967), .A2(new_n984), .A3(new_n771), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n970), .A2(new_n771), .A3(new_n932), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n985), .A2(KEYINPUT53), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(G171), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n975), .A2(new_n982), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(KEYINPUT53), .A3(new_n987), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n980), .A2(G301), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n980), .A2(KEYINPUT127), .A3(G301), .A4(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n991), .B1(new_n974), .B2(G171), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1971), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n969), .A2(new_n1000), .A3(new_n972), .ZN(new_n1001));
  INV_X1    g576(.A(G2090), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n945), .A2(new_n1002), .A3(new_n947), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT55), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1001), .A2(new_n1009), .A3(new_n1003), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1005), .A2(G8), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n930), .B2(new_n933), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT113), .B(G8), .C1(new_n930), .C2(new_n933), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n791), .A2(G1976), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1014), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n605), .B2(KEYINPUT115), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n965), .A2(new_n957), .A3(new_n929), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT113), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1018), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1019), .A2(KEYINPUT116), .A3(new_n1028), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1012), .A2(new_n1021), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n957), .A2(new_n1037), .A3(new_n946), .A4(new_n929), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n947), .A2(KEYINPUT117), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n945), .A2(new_n1038), .A3(new_n1039), .A4(new_n1002), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1001), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1007), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1017), .A2(new_n1018), .B1(G1976), .B2(new_n791), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1012), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1014), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1011), .A2(new_n1036), .A3(new_n1043), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n958), .B2(new_n966), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n945), .A2(new_n742), .A3(new_n947), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G286), .A2(G8), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT123), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT124), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(KEYINPUT51), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1053), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1054), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1052), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1051), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(G286), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n992), .A2(new_n999), .A3(new_n1049), .A4(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1069));
  NOR2_X1   g644(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1070));
  AND2_X1   g645(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1071));
  NOR3_X1   g646(.A1(G299), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n945), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(G2072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n970), .A2(new_n932), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1073), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1029), .A2(G2067), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT120), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n945), .B2(new_n947), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1081), .B1(new_n1085), .B2(new_n621), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1074), .A2(new_n1075), .B1(new_n967), .B2(new_n1078), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1090), .A2(new_n1073), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1029), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n970), .A2(new_n932), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(G1996), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n567), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1099), .A3(new_n567), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1091), .A2(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT61), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1102), .A2(KEYINPUT121), .A3(new_n1080), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1092), .B1(new_n1105), .B2(new_n1076), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1081), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1101), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1101), .B(KEYINPUT122), .C1(new_n1107), .C2(new_n1103), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1085), .A2(KEYINPUT60), .A3(new_n621), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n621), .B1(new_n1085), .B2(KEYINPUT60), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1112), .A2(new_n1113), .B1(KEYINPUT60), .B2(new_n1085), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1068), .B1(new_n1089), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1011), .A2(new_n1036), .A3(new_n1043), .A4(new_n1048), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n989), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1063), .A2(new_n1120), .A3(new_n1066), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1053), .A2(G168), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1036), .A2(new_n1048), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1005), .A2(G8), .A3(new_n1010), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1007), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1124), .A2(new_n1123), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1126), .A2(new_n1011), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1011), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1013), .B1(new_n599), .B2(new_n600), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(G1981), .B2(G305), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1132), .A2(new_n1126), .B1(new_n1136), .B2(new_n1019), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1122), .A2(new_n1131), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n944), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n934), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT48), .Z(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n942), .B2(new_n934), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n934), .B1(new_n938), .B2(new_n726), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n934), .A2(new_n729), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT47), .Z(new_n1149));
  INV_X1    g724(.A(new_n940), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1150), .A2(new_n941), .B1(G2067), .B2(new_n760), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1143), .B(new_n1149), .C1(new_n934), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g728(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1155));
  NOR2_X1   g729(.A1(G229), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n1156), .B(new_n876), .C1(new_n925), .C2(new_n926), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


