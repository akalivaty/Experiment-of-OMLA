//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .A4(G134), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI22_X1  g006(.A1(new_n192), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n192), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n198), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT0), .B(G128), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(new_n202), .B2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(KEYINPUT65), .A3(G143), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n209), .A3(G128), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT0), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n204), .A2(new_n209), .A3(G128), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT67), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n222), .B2(new_n204), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n202), .A2(KEYINPUT65), .A3(G143), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n204), .B2(new_n203), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n216), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n190), .A2(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n192), .A2(G137), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n198), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n188), .A2(new_n189), .B1(new_n190), .B2(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n193), .B2(new_n191), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n231), .B2(new_n198), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n200), .A2(new_n213), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n187), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT0), .A3(G128), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n225), .B2(new_n201), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n197), .B2(new_n199), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n208), .A2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(G128), .B1(new_n215), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n208), .B2(G146), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n206), .B1(new_n243), .B2(new_n240), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n244), .B1(new_n214), .B2(new_n215), .ZN(new_n245));
  INV_X1    g059(.A(new_n229), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n199), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT64), .B(KEYINPUT30), .C1(new_n239), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n235), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G119), .ZN(new_n253));
  INV_X1    g067(.A(G119), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .A3(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(G119), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G113), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(new_n253), .A3(new_n255), .A4(new_n256), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n259), .A2(new_n265), .A3(KEYINPUT69), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT69), .B1(new_n259), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n200), .A2(new_n213), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(new_n265), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n259), .A2(new_n265), .A3(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n226), .A2(new_n232), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n279), .B(KEYINPUT27), .Z(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G101), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n269), .A2(KEYINPUT31), .A3(new_n277), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n268), .B1(new_n239), .B2(new_n248), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT28), .B1(new_n233), .B2(new_n275), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n275), .B1(new_n235), .B2(new_n249), .ZN(new_n293));
  INV_X1    g107(.A(new_n277), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(new_n282), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n284), .B(new_n285), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT32), .B1(new_n296), .B2(G472), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n295), .B2(KEYINPUT31), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n269), .A2(new_n277), .A3(new_n283), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n291), .A3(new_n290), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  INV_X1    g115(.A(G472), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n287), .A2(new_n277), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n305), .B2(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n283), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n293), .A2(new_n294), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n283), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n288), .A2(new_n282), .A3(new_n289), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n311), .B2(KEYINPUT29), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT70), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n316), .B(new_n313), .C1(new_n297), .C2(new_n303), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(G146), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n202), .ZN(new_n324));
  XNOR2_X1  g138(.A(G119), .B(G128), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT71), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n254), .B2(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n254), .A2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G110), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n323), .B(new_n324), .C1(new_n329), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n337), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(G110), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n320), .A2(G146), .A3(new_n322), .ZN(new_n341));
  AOI21_X1  g155(.A(G146), .B1(new_n320), .B2(new_n322), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n325), .B(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n341), .A2(new_n342), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n336), .B(KEYINPUT73), .C1(new_n340), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n335), .B1(new_n344), .B2(new_n327), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n323), .A2(new_n324), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n345), .A2(new_n340), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT22), .B(G137), .ZN(new_n352));
  INV_X1    g166(.A(G953), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n352), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT74), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n336), .B(new_n355), .C1(new_n340), .C2(new_n345), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n359), .B2(KEYINPUT75), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(KEYINPUT75), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n285), .ZN(new_n365));
  INV_X1    g179(.A(new_n362), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n357), .A2(new_n358), .A3(new_n366), .A4(new_n360), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n365), .A2(G902), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT76), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n357), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(KEYINPUT77), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n353), .A2(G227), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT79), .B1(new_n383), .B2(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n383), .A2(KEYINPUT79), .A3(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n394), .A2(new_n392), .A3(G107), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n383), .A2(G104), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n389), .B(new_n393), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n399));
  NOR4_X1   g213(.A1(new_n245), .A2(new_n398), .A3(KEYINPUT81), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n241), .A2(new_n244), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n402), .B2(new_n216), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n388), .A2(new_n397), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT80), .B1(new_n210), .B2(new_n222), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n204), .A2(new_n209), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n202), .A2(G143), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n408), .A2(new_n217), .B1(KEYINPUT1), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n236), .A2(new_n215), .A3(new_n411), .A4(G128), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n399), .B1(new_n413), .B2(new_n398), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n418));
  OAI22_X1  g232(.A1(new_n383), .A2(G104), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n385), .A2(new_n394), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n383), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G104), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n389), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n213), .B(new_n417), .C1(new_n418), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n406), .A2(new_n200), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n200), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n226), .A2(KEYINPUT10), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT81), .B1(new_n428), .B2(new_n398), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n403), .A2(new_n401), .A3(new_n404), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n414), .A2(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n382), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n435));
  INV_X1    g249(.A(new_n382), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n404), .B2(new_n226), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n404), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n245), .A2(new_n398), .A3(KEYINPUT82), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(KEYINPUT12), .A3(new_n200), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT12), .B1(new_n442), .B2(new_n200), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n435), .B(new_n436), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G469), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n285), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n200), .B1(new_n406), .B2(new_n425), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n436), .A3(new_n435), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n200), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n442), .A2(KEYINPUT12), .A3(new_n200), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n427), .ZN(new_n456));
  OAI211_X1 g270(.A(G469), .B(new_n450), .C1(new_n456), .C2(new_n436), .ZN(new_n457));
  NAND2_X1  g271(.A1(G469), .A2(G902), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n448), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n460));
  INV_X1    g274(.A(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n353), .A3(G214), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n208), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n460), .B1(new_n465), .B2(new_n198), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n198), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT86), .A3(G131), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n341), .A2(new_n342), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT86), .B1(new_n469), .B2(G131), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n460), .B(new_n198), .C1(new_n463), .C2(new_n464), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT17), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G113), .B(G122), .Z(new_n477));
  XOR2_X1   g291(.A(KEYINPUT87), .B(G104), .Z(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n465), .B1(new_n480), .B2(new_n198), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(KEYINPUT18), .A3(G131), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n319), .B(new_n202), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n476), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n479), .B1(new_n476), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n285), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT88), .B(G475), .Z(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G478), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G128), .B(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT13), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n208), .A2(G128), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(G134), .C1(KEYINPUT13), .C2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(G116), .B(G122), .Z(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G107), .ZN(new_n498));
  XNOR2_X1  g312(.A(G116), .B(G122), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n383), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n192), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n493), .B(new_n192), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n252), .A2(KEYINPUT14), .A3(G122), .ZN(new_n505));
  OAI211_X1 g319(.A(G107), .B(new_n505), .C1(new_n497), .C2(KEYINPUT14), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT9), .B(G234), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n509), .A2(new_n364), .A3(G953), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n508), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n492), .B1(new_n512), .B2(new_n285), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n508), .A2(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n503), .B2(new_n507), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n285), .B(new_n492), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n319), .B(KEYINPUT19), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n341), .B1(new_n202), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n484), .ZN(new_n524));
  INV_X1    g338(.A(new_n479), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n476), .A2(new_n479), .A3(new_n484), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT20), .B(new_n531), .C1(new_n526), .C2(new_n527), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n489), .B(new_n518), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n353), .A2(G952), .ZN(new_n534));
  INV_X1    g348(.A(G234), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n461), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(G902), .B(G953), .C1(new_n535), .C2(new_n461), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT89), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT21), .B(G898), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G221), .B1(new_n509), .B2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n459), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G210), .B1(G237), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G125), .B1(new_n207), .B2(new_n212), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n226), .B2(G125), .ZN(new_n548));
  INV_X1    g362(.A(G224), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n548), .B(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n252), .A2(G119), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT5), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n260), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n257), .B2(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n404), .A2(new_n265), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G122), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n417), .B1(new_n418), .B2(new_n423), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n558), .C1(new_n275), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT6), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n275), .B2(new_n559), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n552), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n556), .A2(new_n265), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n398), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n558), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n550), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n245), .A2(new_n321), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n547), .ZN(new_n578));
  INV_X1    g392(.A(new_n575), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n548), .A2(new_n579), .B1(KEYINPUT7), .B2(new_n551), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n573), .B(new_n560), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n285), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n546), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n584));
  INV_X1    g398(.A(new_n552), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n560), .A2(KEYINPUT6), .B1(new_n562), .B2(new_n564), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n562), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n569), .A2(new_n398), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n590));
  INV_X1    g404(.A(new_n418), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n415), .A2(G101), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n593), .B2(new_n268), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n594), .A2(new_n558), .B1(new_n571), .B2(new_n572), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n548), .A2(new_n579), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n576), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n548), .A2(new_n574), .A3(KEYINPUT7), .A4(new_n551), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n588), .A2(new_n600), .A3(new_n545), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n583), .A2(new_n584), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G214), .B1(G237), .B2(G902), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT85), .B(new_n546), .C1(new_n568), .C2(new_n582), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n379), .B1(new_n544), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n543), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n457), .A2(new_n458), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n609), .B2(new_n448), .ZN(new_n610));
  INV_X1    g424(.A(new_n605), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT90), .A4(new_n542), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n318), .A2(new_n378), .A3(new_n606), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT91), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  AOI21_X1  g429(.A(new_n545), .B1(new_n588), .B2(new_n600), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n601), .B1(new_n616), .B2(KEYINPUT92), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n618), .B(new_n545), .C1(new_n588), .C2(new_n600), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n603), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT93), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n541), .ZN(new_n623));
  OAI211_X1 g437(.A(KEYINPUT93), .B(new_n603), .C1(new_n617), .C2(new_n619), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n512), .A2(new_n490), .A3(new_n285), .ZN(new_n626));
  NAND2_X1  g440(.A1(G478), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n512), .B(KEYINPUT33), .Z(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(G478), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n489), .B1(new_n530), .B2(new_n532), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n459), .A2(new_n543), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n296), .A2(G472), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n377), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n625), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  OR2_X1    g456(.A1(new_n513), .A2(new_n517), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n643), .B(new_n489), .C1(new_n530), .C2(new_n532), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n625), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT94), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n346), .A2(new_n351), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n346), .B(new_n351), .C1(KEYINPUT36), .C2(new_n356), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n371), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n368), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n638), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n612), .A2(new_n606), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  AND2_X1   g475(.A1(new_n622), .A2(new_n624), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n459), .A2(new_n543), .A3(new_n656), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n537), .B1(new_n539), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n318), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  OAI21_X1  g484(.A(new_n283), .B1(new_n293), .B2(new_n294), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n287), .A2(new_n277), .A3(new_n282), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT97), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(KEYINPUT97), .A3(new_n672), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n285), .A3(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n297), .A2(new_n303), .B1(new_n677), .B2(G472), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n633), .A2(new_n518), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n657), .A3(new_n603), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n665), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n610), .A2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n678), .B(new_n680), .C1(new_n682), .C2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n602), .A2(new_n604), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT96), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n684), .B(new_n686), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n683), .B(new_n688), .C1(KEYINPUT40), .C2(new_n682), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT98), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n208), .ZN(G45));
  NAND2_X1  g505(.A1(new_n634), .A2(new_n666), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n663), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n318), .A2(new_n662), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT99), .B(G146), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G48));
  NAND2_X1  g510(.A1(new_n453), .A2(new_n454), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n382), .B1(new_n455), .B2(new_n427), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n449), .A2(new_n435), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n382), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n543), .A3(new_n448), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n701), .A2(KEYINPUT100), .A3(new_n543), .A4(new_n448), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n704), .A2(new_n634), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n318), .A2(new_n625), .A3(new_n706), .A4(new_n378), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  AND2_X1   g523(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n377), .A2(new_n541), .A3(new_n644), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n318), .A2(new_n662), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT101), .B(G116), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G18));
  AND2_X1   g528(.A1(new_n542), .A2(new_n656), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n318), .A2(new_n662), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  OAI21_X1  g531(.A(KEYINPUT102), .B1(new_n638), .B2(new_n373), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n368), .A2(new_n372), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n637), .A4(new_n636), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n625), .A2(new_n722), .A3(new_n710), .A4(new_n679), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  INV_X1    g538(.A(new_n658), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n692), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n662), .A3(new_n710), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NAND2_X1  g542(.A1(new_n304), .A2(new_n314), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n316), .ZN(new_n730));
  AOI211_X1 g544(.A(G469), .B(G902), .C1(new_n434), .C2(new_n445), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT103), .B1(new_n608), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n603), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n602), .B2(new_n604), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n448), .A2(new_n735), .A3(new_n457), .A4(new_n458), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n543), .A2(new_n732), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n313), .B1(new_n297), .B2(new_n303), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT70), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n730), .A2(new_n737), .A3(new_n739), .A4(new_n378), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n732), .A2(new_n734), .A3(new_n543), .A4(new_n736), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n692), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n729), .B2(new_n719), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n738), .A2(KEYINPUT104), .A3(new_n373), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n741), .A2(new_n742), .B1(new_n748), .B2(KEYINPUT42), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n740), .B2(new_n667), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n315), .A2(new_n317), .A3(new_n377), .ZN(new_n753));
  INV_X1    g567(.A(new_n667), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n754), .A4(new_n737), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  OAI21_X1  g571(.A(new_n450), .B1(new_n456), .B2(new_n436), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n447), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n759), .B2(new_n758), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n458), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n731), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n458), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n607), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n638), .A2(new_n656), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT108), .Z(new_n771));
  AOI21_X1  g585(.A(KEYINPUT43), .B1(new_n633), .B2(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n633), .A2(new_n630), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n633), .B(new_n630), .C1(KEYINPUT107), .C2(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT44), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n734), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n776), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n769), .A2(new_n779), .A3(new_n681), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  XNOR2_X1  g596(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n769), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n769), .B1(KEYINPUT109), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n318), .A2(new_n378), .A3(new_n692), .A4(new_n778), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND2_X1  g603(.A1(new_n701), .A2(new_n448), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT49), .Z(new_n791));
  NOR4_X1   g605(.A1(new_n773), .A2(new_n373), .A3(new_n733), .A4(new_n607), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n687), .A3(new_n678), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n704), .A2(new_n705), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n778), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n536), .B1(new_n774), .B2(new_n775), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n725), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT118), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n796), .A2(new_n722), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n733), .A3(new_n687), .A4(new_n710), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n803));
  AND2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n795), .A2(new_n378), .A3(new_n537), .A4(new_n678), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n632), .A3(new_n630), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n799), .A2(new_n802), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n790), .A2(new_n543), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n784), .B2(new_n786), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n800), .A2(new_n734), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT51), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n807), .B(new_n813), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n797), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n746), .A2(new_n747), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT120), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n800), .A2(new_n662), .A3(new_n710), .ZN(new_n821));
  INV_X1    g635(.A(new_n634), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n821), .B(new_n534), .C1(new_n822), .C2(new_n805), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(KEYINPUT119), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n818), .A2(KEYINPUT120), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT48), .A3(new_n819), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n823), .A2(KEYINPUT119), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT121), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n824), .A2(new_n826), .A3(new_n830), .A4(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n815), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n732), .A2(new_n543), .A3(new_n736), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n656), .A2(new_n665), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n678), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n662), .A4(new_n679), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n677), .A2(G472), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n304), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n607), .B1(new_n459), .B2(KEYINPUT103), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n736), .A3(new_n843), .A4(new_n836), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n622), .A2(new_n624), .A3(new_n679), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n669), .A2(new_n694), .A3(new_n727), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n846), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n622), .A2(new_n624), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n315), .A3(new_n317), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n668), .B2(new_n693), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT52), .A4(new_n727), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT53), .B1(new_n855), .B2(KEYINPUT113), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n756), .A2(new_n749), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n707), .A2(new_n712), .A3(new_n716), .A4(new_n723), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT110), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n644), .B(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n623), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n644), .B(KEYINPUT110), .ZN(new_n864));
  INV_X1    g678(.A(new_n862), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT111), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n639), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n639), .A2(new_n634), .A3(new_n865), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n613), .A2(new_n867), .A3(new_n659), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n533), .A2(new_n665), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT112), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n663), .A3(new_n778), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n318), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n726), .A2(new_n737), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n858), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n855), .A2(new_n857), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n856), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n712), .A2(new_n716), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n707), .A2(new_n723), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT115), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n852), .B(new_n710), .C1(new_n711), .C2(new_n715), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n707), .A4(new_n723), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n613), .A2(new_n867), .A3(new_n659), .A4(new_n868), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n874), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n756), .A3(new_n749), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n881), .A2(new_n877), .B1(new_n892), .B2(new_n855), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n880), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n879), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n880), .A3(new_n894), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n833), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n793), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n353), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n893), .A2(new_n285), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT56), .B1(new_n903), .B2(G210), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n586), .A2(new_n587), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n585), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT122), .B1(new_n893), .B2(new_n285), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n876), .A2(new_n857), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n911), .B2(new_n855), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n849), .A2(new_n854), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n891), .A3(new_n888), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n910), .B(G902), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n909), .A2(new_n915), .A3(new_n546), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n908), .B1(new_n916), .B2(new_n918), .ZN(G51));
  XNOR2_X1  g733(.A(new_n893), .B(KEYINPUT54), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n458), .B(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n446), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n764), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n915), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n901), .B1(new_n922), .B2(new_n924), .ZN(G54));
  AND2_X1   g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n909), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n528), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n902), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n927), .A2(KEYINPUT123), .A3(new_n928), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G60));
  XOR2_X1   g748(.A(new_n629), .B(KEYINPUT124), .Z(new_n935));
  XOR2_X1   g749(.A(new_n627), .B(KEYINPUT59), .Z(new_n936));
  OR2_X1    g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n902), .B1(new_n920), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n936), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n896), .A2(new_n897), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n935), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n893), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n654), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n357), .A2(new_n358), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n893), .B2(new_n943), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n902), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n540), .B2(new_n549), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n858), .A2(new_n869), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n905), .B1(G898), .B2(new_n353), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT125), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n788), .A2(new_n857), .ZN(new_n957));
  INV_X1    g771(.A(new_n848), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n769), .A2(new_n681), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n817), .A2(new_n662), .A3(new_n679), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n781), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n957), .A2(G953), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n664), .A2(new_n353), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G227), .A2(G900), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n250), .B(new_n521), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n964), .A2(G953), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n962), .B2(new_n963), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(G953), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n690), .A2(new_n970), .A3(new_n848), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n690), .B2(new_n848), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n682), .A2(new_n778), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n753), .B(new_n974), .C1(new_n634), .C2(new_n864), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n781), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n973), .A2(new_n788), .A3(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n966), .A2(G953), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n968), .B(new_n969), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n967), .A2(new_n979), .ZN(G72));
  NAND4_X1  g794(.A1(new_n973), .A2(new_n788), .A3(new_n952), .A4(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n671), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n901), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n309), .A2(new_n282), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n878), .A2(new_n671), .A3(new_n988), .A4(new_n983), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(KEYINPUT127), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n957), .A2(new_n961), .A3(new_n858), .A4(new_n869), .ZN(new_n991));
  INV_X1    g805(.A(new_n984), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n987), .A2(new_n989), .A3(new_n993), .ZN(G57));
endmodule


