

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600;

  XOR2_X1 U326 ( .A(n373), .B(n372), .Z(n568) );
  XOR2_X1 U327 ( .A(n315), .B(n451), .Z(n546) );
  NOR2_X2 U328 ( .A1(n496), .A2(n438), .ZN(n439) );
  XNOR2_X2 U329 ( .A(n426), .B(n295), .ZN(n496) );
  XOR2_X2 U330 ( .A(KEYINPUT119), .B(n465), .Z(n580) );
  XOR2_X1 U331 ( .A(KEYINPUT41), .B(n417), .Z(n573) );
  NOR2_X1 U332 ( .A1(n414), .A2(n586), .ZN(n416) );
  XNOR2_X1 U333 ( .A(n380), .B(n379), .ZN(n386) );
  XNOR2_X1 U334 ( .A(n416), .B(n415), .ZN(n425) );
  NOR2_X1 U335 ( .A1(n510), .A2(n593), .ZN(n486) );
  XNOR2_X1 U336 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U337 ( .A(n306), .B(G169GAT), .ZN(n307) );
  XNOR2_X1 U338 ( .A(n491), .B(n490), .ZN(n526) );
  AND2_X1 U339 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U340 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n295) );
  AND2_X1 U341 ( .A1(n482), .A2(n541), .ZN(n296) );
  INV_X1 U342 ( .A(KEYINPUT108), .ZN(n415) );
  XNOR2_X1 U343 ( .A(n378), .B(n294), .ZN(n379) );
  XNOR2_X1 U344 ( .A(n341), .B(n340), .ZN(n380) );
  XOR2_X1 U345 ( .A(n380), .B(n342), .Z(n344) );
  INV_X1 U346 ( .A(KEYINPUT102), .ZN(n485) );
  OR2_X1 U347 ( .A1(n483), .A2(n296), .ZN(n484) );
  XNOR2_X1 U348 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U349 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U350 ( .A(n329), .B(n328), .ZN(n337) );
  NOR2_X1 U351 ( .A1(n546), .A2(n464), .ZN(n465) );
  XNOR2_X1 U352 ( .A(n355), .B(n354), .ZN(n593) );
  INV_X1 U353 ( .A(G134GAT), .ZN(n502) );
  XNOR2_X1 U354 ( .A(KEYINPUT111), .B(n501), .ZN(n556) );
  INV_X1 U355 ( .A(G43GAT), .ZN(n506) );
  XNOR2_X1 U356 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U357 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U358 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U359 ( .A(n505), .B(n504), .ZN(G1343GAT) );
  XNOR2_X1 U360 ( .A(n509), .B(n508), .ZN(G1330GAT) );
  XOR2_X1 U361 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U362 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U363 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U364 ( .A(KEYINPUT19), .B(n299), .ZN(n436) );
  XOR2_X1 U365 ( .A(G190GAT), .B(G134GAT), .Z(n301) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G99GAT), .ZN(n300) );
  XNOR2_X1 U367 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U368 ( .A(G71GAT), .B(KEYINPUT83), .Z(n303) );
  XNOR2_X1 U369 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n302) );
  XNOR2_X1 U370 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U371 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G127GAT), .Z(n342) );
  XOR2_X1 U373 ( .A(n342), .B(G176GAT), .Z(n308) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U376 ( .A(n436), .B(n311), .Z(n315) );
  XOR2_X1 U377 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n313) );
  XNOR2_X1 U378 ( .A(KEYINPUT80), .B(G120GAT), .ZN(n312) );
  XNOR2_X1 U379 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U380 ( .A(G113GAT), .B(n314), .Z(n451) );
  XOR2_X1 U381 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n317) );
  XNOR2_X1 U382 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n317), .B(n316), .ZN(n319) );
  INV_X1 U384 ( .A(KEYINPUT91), .ZN(n318) );
  XNOR2_X1 U385 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U386 ( .A(G148GAT), .B(G78GAT), .Z(n378) );
  XNOR2_X1 U387 ( .A(n378), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n321), .B(n320), .ZN(n323) );
  XNOR2_X1 U389 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n322), .B(KEYINPUT2), .ZN(n446) );
  XOR2_X1 U391 ( .A(n323), .B(n446), .Z(n329) );
  XOR2_X1 U392 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n325) );
  NAND2_X1 U393 ( .A1(G228GAT), .A2(G233GAT), .ZN(n324) );
  XOR2_X1 U394 ( .A(n325), .B(n324), .Z(n327) );
  XOR2_X1 U395 ( .A(G141GAT), .B(G22GAT), .Z(n410) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G162GAT), .Z(n365) );
  XNOR2_X1 U397 ( .A(n410), .B(n365), .ZN(n326) );
  XOR2_X1 U398 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U399 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n333) );
  INV_X1 U401 ( .A(KEYINPUT89), .ZN(n332) );
  XNOR2_X1 U402 ( .A(n333), .B(n332), .ZN(n335) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(G211GAT), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n427) );
  XNOR2_X1 U405 ( .A(n427), .B(KEYINPUT22), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n478) );
  XOR2_X1 U407 ( .A(G64GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U408 ( .A(G211GAT), .B(G155GAT), .ZN(n338) );
  XNOR2_X1 U409 ( .A(n339), .B(n338), .ZN(n355) );
  XOR2_X1 U410 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n341) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G57GAT), .ZN(n340) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U414 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n346) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U417 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U418 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n350) );
  XNOR2_X1 U419 ( .A(G1GAT), .B(G8GAT), .ZN(n349) );
  XNOR2_X1 U420 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n351), .B(KEYINPUT78), .ZN(n352) );
  XNOR2_X1 U422 ( .A(n353), .B(n352), .ZN(n354) );
  INV_X1 U423 ( .A(n593), .ZN(n374) );
  XOR2_X1 U424 ( .A(G134GAT), .B(KEYINPUT76), .Z(n447) );
  XOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .Z(n432) );
  XOR2_X1 U426 ( .A(n447), .B(n432), .Z(n357) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U429 ( .A(G92GAT), .B(KEYINPUT9), .Z(n359) );
  XNOR2_X1 U430 ( .A(KEYINPUT75), .B(KEYINPUT10), .ZN(n358) );
  XNOR2_X1 U431 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U432 ( .A(n361), .B(n360), .Z(n367) );
  XOR2_X1 U433 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n363) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n362) );
  XNOR2_X1 U435 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U436 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n367), .B(n366), .ZN(n373) );
  XOR2_X1 U438 ( .A(G29GAT), .B(G43GAT), .Z(n369) );
  XNOR2_X1 U439 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n369), .B(n368), .ZN(n411) );
  XOR2_X1 U441 ( .A(KEYINPUT71), .B(G85GAT), .Z(n371) );
  XNOR2_X1 U442 ( .A(G99GAT), .B(G106GAT), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n391) );
  XOR2_X1 U444 ( .A(n411), .B(n391), .Z(n372) );
  XOR2_X1 U445 ( .A(KEYINPUT36), .B(n568), .Z(n597) );
  NOR2_X1 U446 ( .A1(n374), .A2(n597), .ZN(n375) );
  XNOR2_X1 U447 ( .A(n375), .B(KEYINPUT45), .ZN(n397) );
  XOR2_X1 U448 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n377) );
  XNOR2_X1 U449 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n377), .B(n376), .ZN(n395) );
  INV_X1 U451 ( .A(n386), .ZN(n384) );
  XOR2_X1 U452 ( .A(KEYINPUT70), .B(KEYINPUT73), .Z(n382) );
  XNOR2_X1 U453 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n381) );
  XOR2_X1 U454 ( .A(n382), .B(n381), .Z(n385) );
  INV_X1 U455 ( .A(n385), .ZN(n383) );
  NAND2_X1 U456 ( .A1(n384), .A2(n383), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n386), .A2(n385), .ZN(n387) );
  NAND2_X1 U458 ( .A1(n388), .A2(n387), .ZN(n393) );
  XOR2_X1 U459 ( .A(G64GAT), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U460 ( .A(G176GAT), .B(G204GAT), .ZN(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n391), .B(n429), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U464 ( .A(n395), .B(n394), .Z(n417) );
  INV_X1 U465 ( .A(n417), .ZN(n396) );
  NAND2_X1 U466 ( .A1(n397), .A2(n396), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n399) );
  NAND2_X1 U468 ( .A1(G229GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U470 ( .A(n400), .B(KEYINPUT29), .Z(n408) );
  XOR2_X1 U471 ( .A(G113GAT), .B(G15GAT), .Z(n402) );
  XNOR2_X1 U472 ( .A(G36GAT), .B(G50GAT), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U474 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n404) );
  XNOR2_X1 U475 ( .A(G197GAT), .B(G1GAT), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U479 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  XOR2_X1 U480 ( .A(n409), .B(n428), .Z(n413) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U482 ( .A(n413), .B(n412), .Z(n528) );
  INV_X1 U483 ( .A(n528), .ZN(n586) );
  NAND2_X1 U484 ( .A1(n586), .A2(n573), .ZN(n418) );
  XNOR2_X1 U485 ( .A(KEYINPUT46), .B(n418), .ZN(n420) );
  NOR2_X1 U486 ( .A1(n593), .A2(n568), .ZN(n419) );
  AND2_X1 U487 ( .A1(n420), .A2(n419), .ZN(n422) );
  INV_X1 U488 ( .A(KEYINPUT47), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n423), .B(KEYINPUT107), .ZN(n424) );
  AND2_X2 U491 ( .A1(n425), .A2(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n435) );
  XNOR2_X1 U493 ( .A(KEYINPUT96), .B(n429), .ZN(n431) );
  NAND2_X1 U494 ( .A1(G226GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n469) );
  BUF_X1 U499 ( .A(n469), .Z(n543) );
  XNOR2_X1 U500 ( .A(n543), .B(KEYINPUT118), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(KEYINPUT54), .ZN(n462) );
  XOR2_X1 U502 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n441) );
  XNOR2_X1 U503 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n443) );
  XNOR2_X1 U506 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U508 ( .A(n445), .B(n444), .Z(n453) );
  XOR2_X1 U509 ( .A(n447), .B(n446), .Z(n449) );
  NAND2_X1 U510 ( .A1(G225GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n461) );
  XOR2_X1 U514 ( .A(G57GAT), .B(G148GAT), .Z(n455) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(G141GAT), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U517 ( .A(G85GAT), .B(G162GAT), .Z(n457) );
  XNOR2_X1 U518 ( .A(G29GAT), .B(G127GAT), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U520 ( .A(n459), .B(n458), .Z(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(n541) );
  NAND2_X1 U522 ( .A1(n462), .A2(n541), .ZN(n584) );
  NOR2_X1 U523 ( .A1(n478), .A2(n584), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT55), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n580), .A2(n568), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n466) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U528 ( .A(n469), .B(KEYINPUT97), .Z(n470) );
  XOR2_X1 U529 ( .A(KEYINPUT27), .B(n470), .Z(n498) );
  INV_X1 U530 ( .A(KEYINPUT28), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n478), .B(n471), .ZN(n549) );
  AND2_X1 U532 ( .A1(n498), .A2(n549), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n546), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n541), .A2(n473), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT98), .ZN(n483) );
  NAND2_X1 U536 ( .A1(n546), .A2(n478), .ZN(n475) );
  XNOR2_X1 U537 ( .A(KEYINPUT26), .B(n475), .ZN(n585) );
  INV_X1 U538 ( .A(n585), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n498), .A2(n476), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n543), .A2(n546), .ZN(n477) );
  NOR2_X1 U541 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n479), .B(KEYINPUT25), .ZN(n480) );
  NAND2_X1 U543 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(n484), .ZN(n510) );
  NOR2_X1 U545 ( .A1(n597), .A2(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n488), .ZN(n540) );
  NOR2_X1 U547 ( .A1(n528), .A2(n417), .ZN(n515) );
  INV_X1 U548 ( .A(n515), .ZN(n489) );
  NOR2_X1 U549 ( .A1(n540), .A2(n489), .ZN(n491) );
  INV_X1 U550 ( .A(KEYINPUT38), .ZN(n490) );
  NOR2_X1 U551 ( .A1(n526), .A2(n541), .ZN(n495) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n493) );
  INV_X1 U553 ( .A(G29GAT), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n541), .A2(n496), .ZN(n497) );
  NAND2_X1 U557 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(KEYINPUT110), .B(n499), .ZN(n561) );
  NOR2_X1 U559 ( .A1(n546), .A2(n561), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n549), .A2(n500), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n556), .A2(n568), .ZN(n505) );
  XOR2_X1 U562 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n503) );
  NOR2_X1 U563 ( .A1(n526), .A2(n546), .ZN(n509) );
  XNOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n507) );
  XOR2_X1 U565 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n513) );
  INV_X1 U566 ( .A(n568), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n593), .A2(n511), .ZN(n512) );
  XNOR2_X1 U568 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n510), .A2(n514), .ZN(n529) );
  NAND2_X1 U570 ( .A1(n515), .A2(n529), .ZN(n523) );
  NOR2_X1 U571 ( .A1(n541), .A2(n523), .ZN(n517) );
  XNOR2_X1 U572 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n516) );
  XNOR2_X1 U573 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U574 ( .A(G1GAT), .B(n518), .Z(G1324GAT) );
  NOR2_X1 U575 ( .A1(n543), .A2(n523), .ZN(n519) );
  XOR2_X1 U576 ( .A(G8GAT), .B(n519), .Z(G1325GAT) );
  NOR2_X1 U577 ( .A1(n546), .A2(n523), .ZN(n521) );
  XNOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U580 ( .A(G15GAT), .B(n522), .Z(G1326GAT) );
  NOR2_X1 U581 ( .A1(n549), .A2(n523), .ZN(n524) );
  XOR2_X1 U582 ( .A(G22GAT), .B(n524), .Z(G1327GAT) );
  NOR2_X1 U583 ( .A1(n526), .A2(n543), .ZN(n525) );
  XOR2_X1 U584 ( .A(G36GAT), .B(n525), .Z(G1329GAT) );
  NOR2_X1 U585 ( .A1(n549), .A2(n526), .ZN(n527) );
  XOR2_X1 U586 ( .A(G50GAT), .B(n527), .Z(G1331GAT) );
  NAND2_X1 U587 ( .A1(n573), .A2(n528), .ZN(n539) );
  INV_X1 U588 ( .A(n539), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n541), .A2(n536), .ZN(n531) );
  XOR2_X1 U591 ( .A(n531), .B(KEYINPUT42), .Z(n532) );
  XNOR2_X1 U592 ( .A(G57GAT), .B(n532), .ZN(G1332GAT) );
  NOR2_X1 U593 ( .A1(n543), .A2(n536), .ZN(n533) );
  XOR2_X1 U594 ( .A(G64GAT), .B(n533), .Z(G1333GAT) );
  NOR2_X1 U595 ( .A1(n546), .A2(n536), .ZN(n535) );
  XNOR2_X1 U596 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(G1334GAT) );
  NOR2_X1 U598 ( .A1(n549), .A2(n536), .ZN(n538) );
  XNOR2_X1 U599 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n538), .B(n537), .ZN(G1335GAT) );
  OR2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n541), .A2(n548), .ZN(n542) );
  XOR2_X1 U603 ( .A(G85GAT), .B(n542), .Z(G1336GAT) );
  NOR2_X1 U604 ( .A1(n543), .A2(n548), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT106), .B(n544), .Z(n545) );
  XNOR2_X1 U606 ( .A(G92GAT), .B(n545), .ZN(G1337GAT) );
  NOR2_X1 U607 ( .A1(n546), .A2(n548), .ZN(n547) );
  XOR2_X1 U608 ( .A(G99GAT), .B(n547), .Z(G1338GAT) );
  NOR2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT44), .B(n550), .Z(n551) );
  XNOR2_X1 U611 ( .A(G106GAT), .B(n551), .ZN(G1339GAT) );
  NAND2_X1 U612 ( .A1(n556), .A2(n586), .ZN(n552) );
  XNOR2_X1 U613 ( .A(n552), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n554) );
  NAND2_X1 U615 ( .A1(n556), .A2(n573), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U617 ( .A(G120GAT), .B(n555), .ZN(G1341GAT) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n558) );
  NAND2_X1 U620 ( .A1(n556), .A2(n593), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n560), .B(n559), .ZN(G1342GAT) );
  NOR2_X1 U623 ( .A1(n585), .A2(n561), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n586), .A2(n569), .ZN(n562) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U627 ( .A1(n569), .A2(n573), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n593), .A2(n569), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT116), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n567), .ZN(G1346GAT) );
  XOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT117), .Z(n571) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n580), .A2(n586), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n580), .A2(n573), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U642 ( .A(G176GAT), .B(KEYINPUT120), .Z(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1349GAT) );
  NAND2_X1 U645 ( .A1(n593), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n590) );
  XOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT124), .Z(n588) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n595) );
  NAND2_X1 U652 ( .A1(n595), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .Z(n592) );
  NAND2_X1 U656 ( .A1(n595), .A2(n417), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1353GAT) );
  NAND2_X1 U658 ( .A1(n593), .A2(n595), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U660 ( .A(n595), .ZN(n596) );
  NOR2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U662 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(G218GAT), .B(n600), .ZN(G1355GAT) );
endmodule

