//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(G57gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT95), .B1(new_n202), .B2(G64gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204));
  INV_X1    g003(.A(G64gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(G57gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n206), .C1(G57gat), .C2(new_n205), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT96), .ZN(new_n208));
  NAND2_X1  g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  OR2_X1    g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n209), .B(new_n210), .C1(new_n214), .C2(new_n211), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT21), .ZN(new_n217));
  NAND2_X1  g016(.A1(G231gat), .A2(G233gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G127gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G1gat), .B2(new_n222), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(G8gat), .Z(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(new_n216), .B2(KEYINPUT21), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n221), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G155gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(G183gat), .B(G211gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n233), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT101), .ZN(new_n237));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT7), .ZN(new_n239));
  NAND2_X1  g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240));
  INV_X1    g039(.A(G85gat), .ZN(new_n241));
  INV_X1    g040(.A(G92gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(KEYINPUT8), .A2(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G99gat), .B(G106gat), .Z(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT97), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n244), .A2(KEYINPUT99), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(KEYINPUT99), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n216), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n245), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(new_n216), .ZN(new_n254));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n251), .B(new_n258), .C1(new_n253), .C2(new_n216), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT100), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(KEYINPUT100), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n257), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n257), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n261), .A2(new_n271), .A3(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n237), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT101), .B(new_n272), .C1(new_n265), .C2(new_n269), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n253), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT17), .ZN(new_n279));
  NOR2_X1   g078(.A1(G29gat), .A2(G36gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT14), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT91), .ZN(new_n283));
  XNOR2_X1  g082(.A(G43gat), .B(G50gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(KEYINPUT15), .B2(new_n284), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G29gat), .ZN(new_n288));
  INV_X1    g087(.A(G36gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT15), .A3(new_n284), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n279), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n287), .A2(new_n279), .A3(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n278), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n291), .ZN(new_n295));
  AND2_X1   g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n253), .A2(new_n295), .B1(KEYINPUT41), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT98), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n298), .B(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n296), .A2(KEYINPUT41), .ZN(new_n303));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n302), .A2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n236), .A2(new_n277), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT102), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n226), .B1(new_n293), .B2(new_n292), .ZN(new_n314));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT92), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n227), .A2(new_n295), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT18), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n314), .A2(KEYINPUT18), .A3(new_n317), .A4(new_n318), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n227), .B(new_n295), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n324));
  XNOR2_X1  g123(.A(new_n316), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G113gat), .B(G141gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G197gat), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT11), .B(G169gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT12), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n332), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n321), .A2(new_n334), .A3(new_n322), .A4(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT36), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340));
  INV_X1    g139(.A(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G113gat), .ZN(new_n342));
  INV_X1    g141(.A(G113gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G120gat), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT1), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G127gat), .A2(G134gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G127gat), .A2(G134gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G134gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n220), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G127gat), .A2(G134gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT68), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n345), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT69), .ZN(new_n355));
  AND2_X1   g154(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n357));
  OAI21_X1  g156(.A(G127gat), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n358), .B(new_n351), .C1(KEYINPUT1), .C2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n354), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n340), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n354), .A2(new_n360), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(KEYINPUT70), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  INV_X1    g167(.A(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(KEYINPUT27), .ZN(new_n371));
  AND2_X1   g170(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n374), .B2(KEYINPUT27), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT27), .B(G183gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n368), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT66), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n371), .ZN(new_n379));
  OR2_X1    g178(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT27), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n369), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT28), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT66), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT26), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n391), .A2(KEYINPUT26), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n369), .A3(new_n381), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(KEYINPUT24), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT24), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G183gat), .A3(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n399), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n391), .B2(KEYINPUT23), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n391), .A2(KEYINPUT23), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n407), .A2(new_n408), .A3(new_n395), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n405), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n407), .A2(new_n411), .A3(new_n408), .A4(new_n395), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n401), .A2(new_n403), .B1(new_n370), .B2(new_n369), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n399), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n363), .A2(new_n367), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n365), .A2(new_n366), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n419), .A2(new_n340), .A3(new_n416), .A4(new_n398), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n425));
  INV_X1    g224(.A(new_n422), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n418), .B2(new_n420), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT73), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n427), .A2(new_n431), .A3(new_n428), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n427), .B2(new_n428), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n420), .A3(new_n426), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT71), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(G15gat), .ZN(new_n441));
  INV_X1    g240(.A(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n436), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT32), .B(new_n435), .C1(new_n445), .C2(new_n437), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n430), .A2(new_n434), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT73), .B1(new_n423), .B2(KEYINPUT34), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n431), .A3(new_n428), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n424), .A3(new_n449), .A4(new_n429), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n446), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n339), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n430), .A2(new_n434), .A3(new_n444), .A4(new_n446), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n451), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT36), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G228gat), .A2(G233gat), .ZN(new_n459));
  AND2_X1   g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT81), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G155gat), .ZN(new_n463));
  INV_X1    g262(.A(G162gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  NAND2_X1  g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(KEYINPUT2), .ZN(new_n470));
  OR2_X1    g269(.A1(G141gat), .A2(G148gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(G141gat), .A2(G148gat), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n475));
  INV_X1    g274(.A(new_n472), .ZN(new_n476));
  NOR2_X1   g275(.A1(G141gat), .A2(G148gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT79), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n471), .A2(new_n479), .A3(new_n472), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n475), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n467), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n474), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G211gat), .B(G218gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G197gat), .B(G204gat), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT74), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(KEYINPUT74), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n487), .A3(new_n491), .A4(new_n489), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n486), .B1(new_n497), .B2(KEYINPUT3), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n459), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n475), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT79), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n479), .B1(new_n471), .B2(new_n472), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n484), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n460), .B1(new_n505), .B2(new_n482), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n504), .A2(new_n506), .B1(new_n469), .B2(new_n473), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT29), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n496), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n498), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  OAI221_X1 g311(.A(new_n498), .B1(new_n499), .B2(new_n459), .C1(new_n509), .C2(new_n510), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(G22gat), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G78gat), .B(G106gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G50gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n513), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT86), .B(G22gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n514), .B(new_n517), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n512), .B2(new_n513), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT87), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n512), .A2(new_n513), .A3(new_n523), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n522), .A2(new_n525), .B1(new_n527), .B2(new_n517), .ZN(new_n528));
  INV_X1    g327(.A(new_n510), .ZN(new_n529));
  NAND2_X1  g328(.A1(G226gat), .A2(G233gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n417), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n530), .B1(new_n398), .B2(new_n416), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G8gat), .B(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(G64gat), .B(G92gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n417), .A2(new_n531), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT29), .B1(new_n398), .B2(new_n416), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(new_n510), .C1(new_n531), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(KEYINPUT77), .A3(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n535), .A2(KEYINPUT30), .A3(new_n541), .A4(new_n538), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n538), .B1(new_n535), .B2(new_n541), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n548), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n486), .A2(KEYINPUT3), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n504), .A2(new_n506), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n508), .A3(new_n474), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n558), .A3(new_n364), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n507), .A4(new_n366), .ZN(new_n560));
  NAND2_X1  g359(.A1(G225gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT4), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n486), .B2(new_n364), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT5), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n486), .A2(new_n364), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n345), .A2(new_n347), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n348), .B1(new_n346), .B2(new_n347), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n351), .A2(KEYINPUT68), .A3(new_n352), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n567), .A2(new_n358), .B1(new_n570), .B2(new_n345), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n557), .A3(new_n474), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n561), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n565), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n571), .B1(new_n486), .B2(KEYINPUT3), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n577), .B2(new_n558), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n365), .A2(new_n562), .A3(new_n507), .A4(new_n366), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(KEYINPUT4), .C1(new_n486), .C2(new_n364), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n572), .B2(KEYINPUT4), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n565), .B(new_n578), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G1gat), .B(G29gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT0), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G85gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT84), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n486), .A2(new_n364), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT82), .B1(new_n596), .B2(new_n562), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n579), .A3(new_n581), .ZN(new_n598));
  AOI211_X1 g397(.A(KEYINPUT5), .B(new_n574), .C1(new_n577), .C2(new_n558), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n598), .A2(new_n599), .B1(new_n564), .B2(new_n575), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n595), .B1(new_n600), .B2(new_n589), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT84), .A3(new_n590), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT6), .B1(new_n600), .B2(new_n589), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n584), .A3(new_n589), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n592), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n594), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n528), .B1(new_n555), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n338), .B1(new_n458), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n517), .B1(new_n520), .B2(new_n526), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n514), .A2(new_n517), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(KEYINPUT87), .B2(new_n524), .ZN(new_n612));
  INV_X1    g411(.A(new_n525), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT83), .B1(new_n605), .B2(new_n592), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT84), .B1(new_n585), .B2(new_n590), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n595), .B(new_n589), .C1(new_n576), .C2(new_n584), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n606), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n593), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n548), .A2(new_n554), .A3(new_n551), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT88), .A3(new_n457), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n559), .B1(new_n582), .B2(new_n583), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n574), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n589), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT39), .B1(new_n573), .B2(new_n574), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n625), .B2(new_n574), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n574), .ZN(new_n632));
  INV_X1    g431(.A(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(KEYINPUT40), .A3(new_n589), .A4(new_n627), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n631), .A2(new_n591), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n614), .B1(new_n621), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n535), .A2(KEYINPUT90), .A3(new_n541), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT37), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640));
  INV_X1    g439(.A(new_n538), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT37), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n535), .A2(KEYINPUT90), .A3(new_n541), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n644), .A2(new_n542), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n605), .A2(new_n592), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n589), .B1(new_n576), .B2(new_n584), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n593), .B1(new_n648), .B2(KEYINPUT89), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT89), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT38), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n645), .A2(new_n649), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n609), .A2(new_n623), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n447), .A2(new_n452), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(new_n555), .A3(new_n607), .A4(new_n528), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT35), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n528), .A2(new_n454), .A3(new_n455), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n621), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT35), .B1(new_n649), .B2(new_n651), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n337), .B1(new_n656), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT94), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT94), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n313), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n620), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n621), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT42), .ZN(new_n673));
  INV_X1    g472(.A(G8gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n668), .B2(new_n621), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT103), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(new_n668), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n679), .B2(new_n457), .ZN(new_n680));
  INV_X1    g479(.A(new_n657), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n679), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n614), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR3_X1   g485(.A1(new_n236), .A2(new_n308), .A3(new_n276), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n666), .B2(new_n667), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n288), .A3(new_n620), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n656), .A2(new_n664), .ZN(new_n694));
  INV_X1    g493(.A(new_n308), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n622), .A2(KEYINPUT104), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n637), .A2(new_n654), .B1(new_n456), .B2(new_n453), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n608), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n664), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n695), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n236), .A2(new_n337), .A3(new_n276), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n607), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n691), .B1(new_n692), .B2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n289), .A3(new_n621), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n555), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  NAND2_X1  g514(.A1(new_n666), .A2(new_n667), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n687), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n442), .B1(new_n717), .B2(new_n681), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n458), .A2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n708), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1330gat));
  AOI21_X1  g521(.A(new_n528), .B1(new_n717), .B2(KEYINPUT107), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n689), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n708), .A2(new_n727), .A3(new_n528), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(G50gat), .B1(new_n723), .B2(new_n725), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT48), .B1(new_n733), .B2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1331gat));
  NAND3_X1  g534(.A1(new_n236), .A2(new_n337), .A3(new_n308), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n277), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n702), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n607), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n202), .ZN(G1332gat));
  AND2_X1   g540(.A1(new_n738), .A2(new_n702), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n555), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n744), .B(new_n745), .Z(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n747), .A3(new_n657), .ZN(new_n748));
  OAI21_X1  g547(.A(G71gat), .B1(new_n739), .B2(new_n457), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n750), .B(new_n751), .Z(G1334gat));
  NAND2_X1  g551(.A1(new_n742), .A2(new_n614), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n236), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n337), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n308), .B1(new_n701), .B2(new_n664), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n658), .A2(KEYINPUT35), .B1(new_n661), .B2(new_n662), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n555), .A2(new_n607), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n699), .B1(new_n761), .B2(new_n614), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT104), .B(new_n528), .C1(new_n555), .C2(new_n607), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(new_n698), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n765), .B2(new_n308), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n759), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n277), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n241), .A3(new_n620), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n277), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n706), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n607), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1336gat));
  OAI21_X1  g574(.A(G92gat), .B1(new_n773), .B2(new_n555), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n276), .A2(new_n242), .A3(new_n621), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT111), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n770), .A2(new_n781), .A3(new_n657), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n773), .B2(new_n457), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n277), .A2(G106gat), .A3(new_n528), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n767), .B2(new_n768), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n614), .B(new_n772), .C1(new_n696), .C2(new_n705), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(KEYINPUT112), .B1(G106gat), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n759), .A2(new_n766), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n759), .A2(new_n766), .A3(KEYINPUT51), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n786), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n789), .A2(G106gat), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n801));
  NAND3_X1  g600(.A1(new_n788), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n785), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n796), .B2(new_n797), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n788), .A2(KEYINPUT112), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n259), .A2(new_n260), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n255), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT100), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n261), .A2(new_n262), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n810), .B2(new_n255), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n259), .A2(new_n256), .A3(new_n260), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n268), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(new_n336), .A3(new_n273), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n819), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n822), .A2(KEYINPUT116), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n271), .B1(new_n812), .B2(new_n813), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n273), .B1(new_n827), .B2(new_n268), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n270), .A2(new_n237), .A3(new_n273), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n323), .A2(new_n325), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n317), .B1(new_n314), .B2(new_n318), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n331), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n335), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n829), .A2(KEYINPUT117), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n276), .B2(new_n834), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n308), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n824), .A2(new_n825), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n820), .A2(new_n273), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n695), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n236), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n736), .A2(new_n276), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n607), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n661), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n336), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n528), .B1(new_n842), .B2(new_n843), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n681), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n607), .A2(new_n621), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT118), .B(new_n528), .C1(new_n842), .C2(new_n843), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n337), .A2(new_n343), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  AOI21_X1  g655(.A(G120gat), .B1(new_n847), .B2(new_n276), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n277), .A2(new_n341), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n854), .B2(new_n858), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n846), .A2(new_n755), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT119), .ZN(new_n861));
  AOI21_X1  g660(.A(G127gat), .B1(new_n860), .B2(KEYINPUT119), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n755), .A2(new_n220), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n861), .A2(new_n862), .B1(new_n854), .B2(new_n863), .ZN(G1342gat));
  NOR3_X1   g663(.A1(new_n308), .A2(new_n357), .A3(new_n356), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n661), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT56), .Z(new_n867));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n695), .A3(new_n852), .A4(new_n853), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT120), .B1(new_n868), .B2(G134gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(G141gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n457), .A2(new_n852), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n614), .A2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n843), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n276), .B2(new_n834), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n829), .A2(new_n877), .A3(new_n830), .A4(new_n834), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n822), .A2(new_n823), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n821), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n308), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n236), .B1(new_n883), .B2(new_n841), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n876), .B1(new_n884), .B2(KEYINPUT122), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n886), .B(new_n236), .C1(new_n883), .C2(new_n841), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n875), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n844), .B2(new_n528), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n873), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n872), .B1(new_n891), .B2(new_n336), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n458), .A2(new_n621), .A3(new_n528), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n845), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G141gat), .A3(new_n337), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n872), .A3(new_n336), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n337), .B(new_n873), .C1(new_n888), .C2(new_n890), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n872), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(G1344gat));
  AND2_X1   g701(.A1(new_n883), .A2(new_n841), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n313), .A2(new_n336), .B1(new_n903), .B2(new_n236), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n614), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n844), .A2(new_n874), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n276), .A2(new_n457), .A3(new_n852), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT59), .B(G148gat), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n910), .A3(new_n276), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n897), .B2(new_n276), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n909), .B(new_n911), .C1(G148gat), .C2(new_n912), .ZN(G1345gat));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n463), .B1(new_n891), .B2(new_n236), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n894), .A2(G155gat), .A3(new_n755), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n463), .A3(new_n236), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n755), .B(new_n873), .C1(new_n888), .C2(new_n890), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n918), .B(KEYINPUT123), .C1(new_n919), .C2(new_n463), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(G1346gat));
  AOI21_X1  g720(.A(new_n464), .B1(new_n891), .B2(new_n695), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n842), .A2(new_n843), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n308), .A2(G162gat), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n620), .A3(new_n893), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n845), .A2(new_n927), .A3(new_n893), .A4(new_n924), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT125), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n928), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  AOI211_X1 g731(.A(new_n308), .B(new_n873), .C1(new_n888), .C2(new_n890), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n931), .B(new_n932), .C1(new_n933), .C2(new_n464), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n620), .A2(new_n555), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n851), .A2(new_n853), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G169gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n337), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n844), .A2(new_n620), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n660), .A2(new_n555), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n336), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n939), .A2(new_n944), .ZN(G1348gat));
  OAI21_X1  g744(.A(G176gat), .B1(new_n937), .B2(new_n277), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n942), .A2(G176gat), .A3(new_n277), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1349gat));
  NAND4_X1  g747(.A1(new_n851), .A2(new_n236), .A3(new_n853), .A4(new_n936), .ZN(new_n949));
  INV_X1    g748(.A(new_n374), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n940), .A2(new_n376), .A3(new_n236), .A4(new_n941), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1350gat));
  AND4_X1   g756(.A1(new_n369), .A2(new_n940), .A3(new_n695), .A4(new_n941), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT126), .ZN(new_n959));
  OAI21_X1  g758(.A(G190gat), .B1(new_n937), .B2(new_n308), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g761(.A(KEYINPUT61), .B(G190gat), .C1(new_n937), .C2(new_n308), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(G1351gat));
  AND2_X1   g763(.A1(new_n936), .A2(new_n457), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n965), .B1(new_n905), .B2(new_n906), .ZN(new_n966));
  OAI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n337), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n458), .A2(new_n555), .A3(new_n528), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n940), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n337), .A2(G197gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR4_X1   g772(.A1(new_n970), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n337), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n277), .A2(G204gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n940), .A2(new_n969), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  OAI21_X1  g777(.A(G204gat), .B1(new_n966), .B2(new_n277), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1353gat));
  OR3_X1    g779(.A1(new_n970), .A2(G211gat), .A3(new_n755), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n236), .B(new_n965), .C1(new_n905), .C2(new_n906), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n966), .B2(new_n308), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n308), .A2(G218gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n970), .B2(new_n987), .ZN(G1355gat));
endmodule


