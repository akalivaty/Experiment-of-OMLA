//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n468), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(new_n469), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n482), .A2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n468), .B2(G114), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(G138), .A3(new_n468), .A4(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n506), .A2(new_n515), .ZN(G166));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n503), .A2(new_n517), .A3(G89), .ZN(new_n518));
  AND3_X1   g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n518), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n518), .A2(new_n529), .A3(new_n522), .A4(new_n526), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n534), .A2(G51), .B1(new_n503), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n528), .A2(new_n530), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  XNOR2_X1  g113(.A(KEYINPUT75), .B(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n503), .A2(new_n517), .A3(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G64), .B1(new_n508), .B2(new_n507), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n505), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n511), .A2(new_n547), .B1(new_n513), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(G56), .B1(new_n508), .B2(new_n507), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n505), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n501), .A2(KEYINPUT78), .A3(new_n502), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n508), .B2(new_n507), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n559), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n511), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n503), .A2(new_n517), .A3(KEYINPUT77), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G91), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT76), .B(KEYINPUT9), .C1(new_n513), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n534), .A2(G53), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n565), .A2(new_n569), .A3(new_n574), .ZN(G299));
  AND2_X1   g150(.A1(new_n543), .A2(new_n544), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n541), .B(new_n540), .C1(new_n576), .C2(new_n505), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  OR2_X1    g153(.A1(new_n503), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n534), .B2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n567), .A2(G87), .A3(new_n568), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n534), .A2(G48), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT80), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n503), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT79), .Z(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n567), .A2(G86), .A3(new_n568), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n505), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n511), .A2(new_n594), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n534), .A2(G54), .ZN(new_n600));
  AND2_X1   g175(.A1(G79), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n560), .A2(new_n562), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n600), .B1(new_n603), .B2(new_n505), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n567), .A2(G92), .A3(new_n568), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .A4(new_n568), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G284));
  XOR2_X1   g185(.A(G284), .B(KEYINPUT81), .Z(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  INV_X1    g192(.A(new_n553), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n612), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n602), .A2(G66), .ZN(new_n620));
  INV_X1    g195(.A(new_n601), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n607), .A2(new_n608), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n467), .A2(new_n465), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n631), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(new_n633), .A3(G2100), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n478), .A2(G2105), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n479), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n468), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n635), .B1(new_n633), .B2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(G2096), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n636), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  NOR2_X1   g244(.A1(G2072), .A2(G2078), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n444), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(KEYINPUT17), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n667), .B(new_n668), .C1(new_n444), .C2(new_n670), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n669), .A3(new_n667), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n683), .A2(new_n688), .A3(new_n686), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n691));
  AOI211_X1 g266(.A(new_n687), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(KEYINPUT103), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1971), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n702), .A2(G23), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G288), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n702), .B1(new_n589), .B2(new_n590), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n702), .A2(G6), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n707), .A2(new_n709), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n711), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n637), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G119), .ZN(new_n723));
  OR2_X1    g298(.A1(G95), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n720), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n702), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n597), .B2(new_n702), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT88), .B(G1986), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n730), .B(new_n734), .C1(KEYINPUT90), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT89), .B1(new_n718), .B2(KEYINPUT34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n718), .A2(KEYINPUT89), .A3(KEYINPUT34), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n735), .A2(KEYINPUT90), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT91), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n737), .B(new_n743), .C1(new_n738), .C2(new_n740), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n720), .A2(G35), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT101), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n720), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n752), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G168), .A2(new_n702), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n702), .B2(G21), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n720), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n720), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(new_n443), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n467), .A2(G141), .A3(new_n468), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n467), .A2(G129), .A3(G2105), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n465), .A2(G105), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n766), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G29), .B2(G32), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n758), .A2(new_n759), .B1(new_n776), .B2(new_n775), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n761), .A2(new_n764), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G116), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n464), .B1(new_n781), .B2(G2105), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT95), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n467), .A2(G140), .A3(new_n468), .ZN(new_n791));
  OAI211_X1 g366(.A(G128), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT96), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n720), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n702), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  INV_X1    g377(.A(G299), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n702), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1956), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n780), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n702), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n609), .B2(new_n702), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT92), .B(G1348), .Z(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G171), .A2(new_n702), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G5), .B2(new_n702), .ZN(new_n814));
  INV_X1    g389(.A(G1961), .ZN(new_n815));
  INV_X1    g390(.A(G2084), .ZN(new_n816));
  AND2_X1   g391(.A1(KEYINPUT24), .A2(G34), .ZN(new_n817));
  NOR2_X1   g392(.A1(KEYINPUT24), .A2(G34), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n720), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  INV_X1    g395(.A(G160), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n720), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n814), .A2(new_n815), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n816), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n720), .A2(G33), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n467), .A2(G139), .A3(new_n468), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT97), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n468), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n829), .A2(KEYINPUT98), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n828), .B(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n827), .B1(new_n841), .B2(new_n720), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(G2072), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(G2072), .ZN(new_n844));
  INV_X1    g419(.A(G28), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT30), .ZN(new_n846));
  AOI21_X1  g421(.A(G29), .B1(new_n845), .B2(KEYINPUT30), .ZN(new_n847));
  OR2_X1    g422(.A1(KEYINPUT31), .A2(G11), .ZN(new_n848));
  NAND2_X1  g423(.A1(KEYINPUT31), .A2(G11), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n846), .A2(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n644), .B2(new_n720), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n702), .A2(G19), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n553), .B2(new_n702), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1341), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n826), .A2(new_n843), .A3(new_n844), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n810), .B2(new_n811), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n807), .A2(new_n812), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n701), .B1(new_n747), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g435(.A(KEYINPUT103), .B(new_n858), .C1(new_n745), .C2(new_n746), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(G311));
  NAND2_X1  g437(.A1(new_n747), .A2(new_n859), .ZN(G150));
  NOR2_X1   g438(.A1(new_n625), .A2(new_n616), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n503), .A2(G67), .ZN(new_n866));
  AND2_X1   g441(.A1(G80), .A2(G543), .ZN(new_n867));
  OAI21_X1  g442(.A(G651), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n503), .A2(new_n517), .A3(G93), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  OAI211_X1 g445(.A(G55), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n618), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n553), .B(new_n868), .C1(new_n873), .C2(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n865), .B(new_n877), .Z(new_n878));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n879));
  AOI21_X1  g454(.A(G860), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n879), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT105), .ZN(G145));
  NAND2_X1  g460(.A1(new_n791), .A2(new_n792), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n787), .B2(new_n789), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n499), .A2(new_n497), .ZN(new_n888));
  INV_X1    g463(.A(new_n495), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n887), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n773), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n772), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n793), .A2(G164), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n887), .A2(new_n890), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n841), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n772), .B1(new_n891), .B2(new_n892), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n837), .A2(new_n839), .ZN(new_n901));
  INV_X1    g476(.A(new_n772), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n637), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n479), .A2(G130), .ZN(new_n906));
  OR2_X1    g481(.A1(G106), .A2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n899), .B2(new_n904), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n911), .A2(new_n630), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n899), .A2(new_n904), .ZN(new_n914));
  INV_X1    g489(.A(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n631), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n726), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n630), .B1(new_n911), .B2(new_n912), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n631), .A3(new_n910), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n727), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n644), .A2(G160), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n644), .A2(G160), .ZN(new_n923));
  INV_X1    g498(.A(G162), .ZN(new_n924));
  OR3_X1    g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n918), .A2(new_n921), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n918), .A2(new_n933), .A3(new_n930), .A4(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n918), .A2(new_n921), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n925), .A2(new_n927), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n935), .A2(KEYINPUT40), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT40), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(G395));
  XNOR2_X1  g516(.A(new_n877), .B(KEYINPUT108), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(new_n626), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n625), .A2(new_n803), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n623), .A2(new_n624), .A3(G299), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n609), .B2(G299), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n625), .A2(KEYINPUT109), .A3(new_n803), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT41), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n609), .B2(G299), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n944), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI221_X1 g533(.A(new_n947), .B1(KEYINPUT110), .B2(new_n956), .C1(new_n943), .C2(new_n954), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n589), .A2(new_n590), .A3(G290), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G290), .B1(new_n589), .B2(new_n590), .ZN(new_n962));
  INV_X1    g537(.A(G288), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(G303), .ZN(new_n964));
  NOR2_X1   g539(.A1(G288), .A2(G166), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n961), .A2(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n962), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n960), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(KEYINPUT110), .B2(new_n956), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n958), .A2(new_n959), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n958), .B2(new_n959), .ZN(new_n974));
  OAI21_X1  g549(.A(G868), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n874), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(G868), .B2(new_n976), .ZN(G295));
  OAI21_X1  g552(.A(new_n975), .B1(G868), .B2(new_n976), .ZN(G331));
  NAND2_X1  g553(.A1(new_n530), .A2(new_n536), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n522), .A2(new_n526), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n529), .B1(new_n980), .B2(new_n518), .ZN(new_n981));
  OAI21_X1  g556(.A(G301), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(G171), .A2(new_n528), .A3(new_n530), .A4(new_n536), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n875), .A2(new_n876), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT112), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n875), .A2(new_n876), .B1(new_n982), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n983), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n877), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n946), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n877), .A2(new_n989), .A3(KEYINPUT111), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n877), .A2(new_n989), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT111), .A3(new_n984), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n991), .B(new_n970), .C1(new_n954), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n954), .B2(new_n995), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n970), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n991), .B(KEYINPUT113), .C1(new_n954), .C2(new_n995), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT41), .B1(new_n944), .B2(new_n945), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n990), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n993), .A2(KEYINPUT112), .A3(new_n984), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n995), .A2(new_n946), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n970), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT43), .B1(new_n1018), .B2(new_n998), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n999), .A2(new_n1000), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n971), .A3(new_n1002), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n996), .A2(new_n997), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1004), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1018), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1021), .B(new_n1022), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n949), .A2(new_n950), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(new_n953), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1014), .B1(new_n1031), .B2(new_n1008), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1017), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n971), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1004), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1021), .B1(new_n1036), .B2(new_n1022), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1020), .B1(new_n1029), .B2(new_n1037), .ZN(G397));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n890), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT116), .B(KEYINPUT45), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G160), .A2(G40), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n793), .A2(G2067), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n887), .A2(new_n799), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1048), .B2(new_n772), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1044), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n1050), .B2(G1996), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  INV_X1    g627(.A(G1996), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1044), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(KEYINPUT46), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(KEYINPUT46), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1049), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n895), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n772), .A2(G1996), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1050), .B1(new_n1047), .B2(new_n1061), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1060), .A2(KEYINPUT118), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT118), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n727), .A2(new_n729), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n727), .A2(new_n729), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1044), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT127), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1063), .A2(KEYINPUT127), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1050), .A2(G1986), .A3(G290), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1072), .B(KEYINPUT48), .Z(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1046), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1044), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1059), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n584), .A2(new_n1079), .A3(new_n590), .A4(new_n588), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n503), .A2(new_n517), .A3(G86), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n584), .A2(new_n588), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G1981), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G164), .A2(G1384), .ZN(new_n1087));
  INV_X1    g662(.A(G40), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n471), .A2(new_n474), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT49), .B1(new_n1084), .B2(new_n1080), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1090), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1089), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1040), .A2(KEYINPUT50), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT119), .B(G2090), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1087), .A2(KEYINPUT45), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1042), .A3(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(G1971), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(G166), .B2(new_n1086), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1107), .A2(new_n1113), .A3(G8), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n963), .A2(G1976), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1090), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT52), .ZN(new_n1118));
  INV_X1    g693(.A(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(G288), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1090), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1118), .B(new_n1121), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1095), .A2(new_n1096), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1041), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1043), .B1(new_n1087), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT45), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1040), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1966), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1098), .A2(new_n1099), .A3(G2084), .ZN(new_n1130));
  OAI21_X1  g705(.A(G8), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G286), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1100), .A2(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1111), .B1(new_n1133), .B2(new_n1086), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1115), .A2(new_n1124), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1107), .A2(G8), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1122), .B1(new_n1138), .B2(new_n1111), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(KEYINPUT63), .A3(new_n1115), .A4(new_n1132), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1123), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1103), .A2(new_n1042), .A3(new_n1089), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1100), .B2(G1956), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n565), .A2(KEYINPUT121), .A3(new_n569), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n1146));
  AND3_X1   g721(.A1(G299), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G299), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g725(.A(new_n1143), .B1(new_n1148), .B2(new_n1147), .C1(new_n1100), .C2(G1956), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1043), .B1(KEYINPUT50), .B2(new_n1040), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1348), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n609), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1150), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1150), .A2(KEYINPUT61), .A3(new_n1151), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  OAI221_X1 g737(.A(new_n625), .B1(G2067), .B2(new_n1156), .C1(new_n1100), .C2(G1348), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n1158), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1160), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1104), .B2(G1996), .ZN(new_n1168));
  AND4_X1   g743(.A1(KEYINPUT122), .A2(new_n1168), .A3(KEYINPUT59), .A4(new_n553), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1168), .B2(new_n553), .ZN(new_n1171));
  NOR4_X1   g746(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n625), .A4(new_n1157), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1159), .B1(new_n1165), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1115), .A2(new_n1124), .A3(new_n1134), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1103), .A2(new_n1042), .A3(new_n443), .A4(new_n1089), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n815), .A2(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1126), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1128), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G171), .B(KEYINPUT54), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1042), .A2(new_n1089), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1184), .A2(KEYINPUT124), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(KEYINPUT124), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n443), .A2(KEYINPUT125), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1178), .B1(KEYINPUT125), .B2(new_n443), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1103), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1190), .A2(new_n1179), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1183), .B1(new_n1191), .B2(new_n1182), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n759), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1153), .A2(new_n816), .A3(new_n1154), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1194), .A2(KEYINPUT123), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1196), .A2(new_n1198), .A3(G168), .ZN(new_n1199));
  AND2_X1   g774(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1200));
  NOR2_X1   g775(.A1(G168), .A2(new_n1086), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1201), .A2(KEYINPUT51), .ZN(new_n1202));
  AOI22_X1  g777(.A1(new_n1199), .A2(new_n1200), .B1(new_n1131), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1201), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1175), .B(new_n1192), .C1(new_n1203), .C2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1141), .B1(new_n1174), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(G301), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1139), .A2(new_n1115), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1131), .A2(new_n1202), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1205), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1209), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1214), .A2(KEYINPUT126), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1216), .B1(new_n1214), .B2(KEYINPUT126), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1207), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1068), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n597), .B(G1986), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1219), .B1(new_n1050), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1078), .B1(new_n1218), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g797(.A1(G227), .A2(new_n462), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n699), .A2(new_n665), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n935), .A2(new_n938), .ZN(new_n1226));
  AND3_X1   g800(.A1(new_n1225), .A2(new_n1226), .A3(new_n1036), .ZN(G308));
  NAND3_X1  g801(.A1(new_n1225), .A2(new_n1226), .A3(new_n1036), .ZN(G225));
endmodule


