//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT66), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n469), .A3(G125), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n476), .A2(new_n469), .A3(KEYINPUT64), .A4(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n473), .A2(new_n475), .B1(G2105), .B2(new_n482), .ZN(G160));
  NAND4_X1  g058(.A1(new_n465), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n470), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT68), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n468), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AND4_X1   g075(.A1(G2105), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G126), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n476), .A2(new_n469), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n502), .A2(new_n510), .A3(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n505), .A2(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  INV_X1    g088(.A(new_n495), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n498), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT69), .B1(new_n498), .B2(G2105), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G126), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n484), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n512), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n528), .A2(G651), .B1(new_n532), .B2(G50), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n529), .A2(new_n530), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n524), .A2(new_n525), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n538), .B(KEYINPUT71), .C1(new_n530), .C2(new_n529), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n533), .B1(new_n534), .B2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT7), .Z(new_n544));
  NAND3_X1  g119(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n544), .B(new_n546), .C1(G51), .C2(new_n532), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n537), .A2(new_n539), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G89), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n548), .A2(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n526), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(new_n532), .B2(G52), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND2_X1  g132(.A1(new_n548), .A2(G81), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G651), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n561), .A2(new_n562), .B1(G43), .B2(new_n532), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT72), .B1(new_n559), .B2(new_n560), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n558), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G860), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT73), .ZN(G188));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n531), .A2(KEYINPUT74), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT74), .B1(new_n531), .B2(new_n573), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n538), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n560), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n537), .A2(G91), .A3(new_n539), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT75), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  OAI21_X1  g158(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT76), .Z(new_n585));
  NAND2_X1  g160(.A1(new_n548), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n532), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n532), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n524), .B2(new_n525), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n537), .A2(G86), .A3(new_n539), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n526), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n532), .B2(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n540), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n548), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n540), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n538), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n613), .A2(new_n560), .B1(new_n614), .B2(new_n531), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n607), .B1(new_n616), .B2(G868), .ZN(G284));
  XNOR2_X1  g192(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G168), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT80), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n581), .B(KEYINPUT75), .Z(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n622), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(G868), .B2(new_n622), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n565), .A2(new_n619), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n612), .A2(new_n615), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n507), .A2(new_n462), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n637));
  INV_X1    g212(.A(G123), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n484), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n491), .B2(G135), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT83), .ZN(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n665), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n684), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT87), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n682), .A2(new_n688), .A3(new_n684), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G24), .B(G290), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1986), .Z(new_n702));
  NOR2_X1   g277(.A1(G25), .A2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n468), .A2(G107), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n484), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n491), .B2(G131), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(G29), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n702), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT89), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1971), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(G23), .ZN(new_n719));
  INV_X1    g294(.A(G288), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n714), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G6), .B(G305), .S(G16), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n718), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n713), .B1(new_n727), .B2(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(G168), .A2(G16), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(KEYINPUT98), .C1(G16), .C2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT98), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G26), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT91), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g318(.A(G128), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n468), .A2(G116), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n484), .A2(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n491), .B2(G140), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n743), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n714), .A2(G4), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n616), .B2(new_n714), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n752), .B1(G1348), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n641), .A2(new_n740), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT30), .B(G28), .Z(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n714), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n714), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n756), .B(new_n759), .C1(new_n761), .C2(G1961), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n762), .B1(G1348), .B2(new_n754), .C1(G1961), .C2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(G160), .A2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(KEYINPUT24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT24), .B2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G2084), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n714), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n565), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n740), .A2(G32), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT26), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n777), .A2(new_n778), .B1(G105), .B2(new_n462), .ZN(new_n779));
  INV_X1    g354(.A(G129), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n484), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G141), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n470), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n774), .B1(new_n785), .B2(new_n740), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n773), .A2(G1341), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G1341), .B2(new_n773), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n763), .A2(new_n770), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n755), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT100), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n622), .B2(new_n714), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n740), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n740), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G2078), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G2078), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n798), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G29), .A2(G35), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G162), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT29), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G2090), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(G2090), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n792), .A2(new_n805), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n491), .A2(G139), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n507), .A2(G127), .ZN(new_n818));
  INV_X1    g393(.A(G115), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n461), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n813), .B(new_n817), .C1(G2105), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  NOR2_X1   g397(.A1(G29), .A2(G33), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT92), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  INV_X1    g401(.A(G2072), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT96), .ZN(new_n829));
  INV_X1    g404(.A(new_n786), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n830), .A2(new_n787), .B1(G2084), .B2(new_n769), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n826), .A2(new_n827), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n826), .A2(KEYINPUT95), .A3(new_n827), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT97), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n829), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT101), .B1(new_n812), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n755), .A2(new_n811), .A3(new_n791), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n804), .A3(new_n809), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n845), .A2(new_n846), .A3(new_n841), .A4(new_n839), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n733), .A2(new_n734), .B1(new_n843), .B2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n734), .A2(new_n733), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(G150));
  NAND2_X1  g426(.A1(new_n616), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n532), .A2(G55), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n854), .B1(new_n560), .B2(new_n855), .C1(new_n540), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n565), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n565), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n853), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n566), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(G145));
  NOR2_X1   g443(.A1(new_n513), .A2(new_n519), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n748), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n821), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n784), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n708), .B(new_n633), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n491), .A2(G142), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT103), .Z(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G118), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(G2105), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n501), .B2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n873), .B(new_n880), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n641), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n881), .B(KEYINPUT104), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n872), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n884), .B1(new_n882), .B2(new_n886), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g467(.A1(new_n857), .A2(new_n619), .ZN(new_n893));
  XNOR2_X1  g468(.A(G288), .B(G305), .ZN(new_n894));
  XOR2_X1   g469(.A(G303), .B(G290), .Z(new_n895));
  XOR2_X1   g470(.A(new_n894), .B(new_n895), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT42), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n622), .A2(new_n628), .A3(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n622), .A2(new_n628), .ZN(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n616), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT41), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n629), .B(new_n860), .ZN(new_n910));
  MUX2_X1   g485(.A(new_n904), .B(new_n909), .S(new_n910), .Z(new_n911));
  OR2_X1    g486(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n911), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n912), .A2(new_n913), .B1(new_n898), .B2(new_n897), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n893), .B1(new_n914), .B2(new_n619), .ZN(G295));
  NAND2_X1  g490(.A1(G295), .A2(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(new_n893), .C1(new_n914), .C2(new_n619), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  AOI21_X1  g495(.A(G168), .B1(new_n920), .B2(G301), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(G301), .A2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n858), .A2(new_n924), .A3(new_n859), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n858), .B2(new_n859), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n860), .A2(new_n923), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n921), .A3(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n905), .A3(new_n908), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n900), .A3(new_n903), .A4(new_n930), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n896), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n888), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n896), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n936), .A3(new_n933), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n926), .A2(new_n927), .A3(new_n922), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n921), .B1(new_n929), .B2(new_n925), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n942), .A2(new_n943), .B1(new_n907), .B2(new_n906), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT41), .B1(new_n900), .B2(new_n903), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n906), .A2(new_n907), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n931), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n950), .A3(new_n933), .ZN(new_n951));
  INV_X1    g526(.A(new_n896), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n935), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(KEYINPUT43), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n941), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n940), .B2(new_n957), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g536(.A(KEYINPUT125), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(new_n965), .C1(new_n513), .C2(new_n519), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n473), .A2(new_n475), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n482), .A2(G2105), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n967), .A3(G40), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT115), .B(G2084), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n511), .B2(new_n520), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n970), .B(new_n971), .C1(new_n964), .C2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n965), .B1(new_n513), .B2(new_n519), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(G160), .A3(G40), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n511), .B2(new_n520), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n738), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n963), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT114), .B(G8), .Z(new_n983));
  NOR2_X1   g558(.A1(G168), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT51), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(KEYINPUT51), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT70), .B1(new_n502), .B2(new_n510), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n513), .A2(new_n519), .A3(new_n512), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n965), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n969), .B1(new_n989), .B2(KEYINPUT50), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n521), .A2(new_n978), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  AOI221_X4 g567(.A(new_n992), .B1(new_n482), .B2(G2105), .C1(new_n473), .C2(new_n475), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n993), .A3(new_n976), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n990), .A2(new_n971), .B1(new_n994), .B2(new_n738), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(new_n995), .B2(new_n983), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n985), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT62), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n999));
  INV_X1    g574(.A(new_n984), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n973), .A2(new_n981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n984), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n997), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n993), .B(new_n966), .C1(new_n972), .C2(new_n964), .ZN(new_n1006));
  INV_X1    g581(.A(G1961), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n977), .A2(G2078), .A3(new_n980), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(KEYINPUT123), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n991), .A2(new_n1013), .A3(new_n993), .A4(new_n976), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n978), .B1(new_n513), .B2(new_n519), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n967), .A2(new_n1018), .A3(G40), .A4(new_n968), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n989), .B2(new_n975), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT53), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT55), .ZN(new_n1025));
  AOI211_X1 g600(.A(KEYINPUT50), .B(G1384), .C1(new_n511), .C2(new_n520), .ZN(new_n1026));
  INV_X1    g601(.A(new_n974), .ZN(new_n1027));
  OAI211_X1 g602(.A(G160), .B(G40), .C1(new_n1027), .C2(new_n964), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2090), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n993), .B(new_n1018), .C1(new_n972), .C2(KEYINPUT45), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1025), .B1(new_n1033), .B2(new_n983), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1020), .B2(G1971), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(KEYINPUT113), .A3(new_n1032), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n990), .A2(new_n1030), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1025), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n993), .A2(new_n1027), .ZN(new_n1042));
  INV_X1    g617(.A(new_n983), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(new_n1043), .C1(new_n1044), .C2(G288), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n967), .A2(G40), .A3(new_n968), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n974), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n983), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n597), .A2(new_n1050), .A3(new_n598), .A4(new_n599), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n599), .A2(new_n598), .ZN(new_n1052));
  OAI21_X1  g627(.A(G1981), .B1(new_n1052), .B2(new_n596), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1053), .A3(KEYINPUT49), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1049), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n720), .A2(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1049), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1046), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1023), .A2(new_n1034), .A3(new_n1041), .A4(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n962), .B1(new_n1005), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n985), .A2(new_n996), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(new_n998), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1041), .A2(new_n1034), .A3(new_n1062), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n976), .A2(G40), .A3(G160), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT123), .A3(new_n1013), .A4(new_n991), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1008), .ZN(new_n1071));
  OAI21_X1  g646(.A(G171), .B1(new_n1071), .B2(new_n1021), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1065), .A2(new_n998), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT125), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1064), .A2(new_n1066), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1046), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n521), .B2(new_n965), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1032), .B1(new_n1078), .B2(new_n1019), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1079), .A2(new_n1035), .B1(new_n990), .B2(new_n1030), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n963), .B1(new_n1080), .B2(new_n1037), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1081), .B2(new_n1040), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n995), .A2(G286), .A3(new_n983), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1034), .A4(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1041), .A2(new_n1034), .A3(new_n1062), .A4(new_n1084), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT116), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1039), .A2(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1091), .B2(new_n1025), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1092), .A2(new_n1082), .A3(KEYINPUT118), .A4(new_n1084), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1089), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1019), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1013), .C1(KEYINPUT45), .C2(new_n972), .ZN(new_n1099));
  AOI21_X1  g674(.A(G171), .B1(new_n1099), .B2(new_n1010), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1070), .A2(new_n1008), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1047), .A2(KEYINPUT124), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NAND3_X1  g678(.A1(G160), .A2(new_n1103), .A3(G40), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1018), .A2(KEYINPUT53), .A3(new_n1013), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1102), .A2(new_n1104), .A3(new_n976), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1008), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G171), .B1(new_n1107), .B2(new_n1021), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1101), .A2(KEYINPUT54), .A3(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1065), .A2(new_n1109), .A3(new_n1067), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1107), .A2(new_n1021), .A3(G171), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1023), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT56), .B(G2072), .Z(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n1031), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n797), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n989), .A2(new_n975), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1114), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1098), .A4(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n581), .B(KEYINPUT57), .Z(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1115), .A2(KEYINPUT120), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n964), .B1(new_n521), .B2(new_n965), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n969), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1047), .A2(G2067), .A3(new_n974), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1131), .A2(new_n628), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n628), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT60), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1098), .B(new_n1137), .C1(KEYINPUT45), .C2(new_n972), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1042), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n565), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(KEYINPUT121), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n628), .A2(KEYINPUT60), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1132), .B1(new_n1006), .B2(new_n1129), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1141), .A2(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1136), .A2(new_n1143), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1121), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1124), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT61), .B1(new_n1151), .B2(new_n1122), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1128), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1135), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1122), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1110), .B(new_n1113), .C1(new_n1153), .C2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1041), .A2(new_n1077), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1058), .A2(new_n1044), .A3(new_n720), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1051), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1049), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1076), .A2(new_n1097), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1047), .A2(new_n976), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1137), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT111), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1163), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n748), .B(G2067), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(G1996), .B2(new_n784), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1165), .A2(new_n784), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT112), .Z(new_n1171));
  AND2_X1   g746(.A1(new_n708), .A2(new_n710), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n708), .A2(new_n710), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1163), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(G290), .B(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1163), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1165), .B(KEYINPUT46), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1163), .B1(new_n1168), .B2(new_n784), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1175), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n748), .A2(new_n750), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1166), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1178), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1178), .A2(KEYINPUT126), .A3(new_n1189), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n459), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n699), .A2(new_n663), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n891), .A2(new_n1198), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n959), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1196), .B1(new_n959), .B2(new_n1199), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n1201), .ZN(G308));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n1199), .ZN(G225));
endmodule


