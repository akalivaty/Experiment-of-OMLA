//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(KEYINPUT67), .A3(G101), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT68), .ZN(G160));
  INV_X1    g051(.A(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n462), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n485), .A2(new_n462), .A3(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n485), .B2(new_n462), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(new_n494), .B2(G114), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n482), .A2(new_n503), .A3(G138), .A4(new_n462), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT71), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(new_n506), .A3(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(G543), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  AND2_X1   g097(.A1(new_n516), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n512), .A2(G89), .A3(new_n516), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n531), .A3(new_n526), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT72), .B1(new_n533), .B2(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n514), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G52), .Z(new_n539));
  OAI22_X1  g114(.A1(new_n517), .A2(new_n538), .B1(new_n520), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT74), .B(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n517), .A2(new_n544), .B1(new_n520), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT75), .B1(new_n543), .B2(new_n546), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n520), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n523), .A2(new_n560), .A3(G53), .ZN(new_n561));
  INV_X1    g136(.A(new_n517), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n559), .A2(new_n561), .B1(new_n562), .B2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n512), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(KEYINPUT76), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n523), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n512), .A2(G87), .A3(new_n516), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n523), .A2(G48), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n514), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n512), .A2(G86), .A3(new_n516), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  XOR2_X1   g157(.A(KEYINPUT77), .B(G85), .Z(new_n583));
  AOI22_X1  g158(.A1(new_n562), .A2(new_n583), .B1(G47), .B2(new_n523), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n514), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  OR3_X1    g165(.A1(G171), .A2(KEYINPUT78), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(G171), .B2(new_n590), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n562), .A2(KEYINPUT10), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n509), .A2(new_n511), .ZN(new_n599));
  INV_X1    g174(.A(new_n507), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n591), .B(new_n592), .C1(G868), .C2(new_n606), .ZN(G284));
  XOR2_X1   g182(.A(G284), .B(KEYINPUT79), .Z(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n606), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g191(.A1(new_n467), .A2(new_n468), .ZN(new_n617));
  INV_X1    g192(.A(new_n460), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT13), .Z(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n479), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n627), .C1(new_n628), .C2(new_n483), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n621), .B2(new_n622), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n649), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n662), .A2(new_n663), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n667), .A2(KEYINPUT82), .A3(new_n668), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n686));
  AND2_X1   g261(.A1(G288), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT87), .A4(new_n575), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n690), .B2(new_n684), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(KEYINPUT33), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(KEYINPUT33), .ZN(new_n693));
  AOI21_X1  g268(.A(G1976), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G22), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G166), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n698), .A2(G1971), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(G1971), .B1(new_n698), .B2(new_n699), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n694), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n692), .A2(G1976), .A3(new_n693), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n684), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n581), .B2(new_n684), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(KEYINPUT86), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(KEYINPUT86), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  NAND3_X1  g285(.A1(new_n702), .A2(new_n703), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n702), .A2(new_n713), .A3(new_n710), .A4(new_n703), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n617), .A2(G2105), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n479), .A2(G119), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n462), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT85), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT84), .B(G29), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G25), .B2(new_n723), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G24), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n588), .B2(G16), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n712), .A2(new_n714), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n722), .A2(G35), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT96), .Z(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n722), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n723), .A2(G27), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n723), .ZN(new_n742));
  INV_X1    g317(.A(G2078), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n684), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n684), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n740), .B(new_n744), .C1(G1961), .C2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n715), .A2(G141), .B1(new_n479), .B2(G129), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n460), .A2(G105), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n722), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n715), .A2(G140), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n479), .A2(G128), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(new_n755), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n757), .A2(new_n758), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT31), .B(G11), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n629), .A2(new_n722), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n759), .A2(new_n770), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n746), .A2(G1961), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n739), .B2(G2090), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n747), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n755), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n482), .A2(G139), .A3(new_n462), .ZN(new_n787));
  AOI21_X1  g362(.A(KEYINPUT90), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(KEYINPUT90), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  INV_X1    g366(.A(G127), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n617), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n482), .A2(G127), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n462), .B1(new_n797), .B2(new_n791), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n789), .A2(new_n790), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n783), .B1(new_n800), .B2(new_n755), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(G160), .A2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n722), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G2084), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n684), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n684), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n802), .B(new_n809), .C1(G1966), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n684), .A2(G20), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT23), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G299), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G1956), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n811), .A2(KEYINPUT95), .A3(G1966), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT95), .B1(new_n811), .B2(G1966), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n782), .A2(new_n812), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n552), .A2(new_n684), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n684), .B2(G19), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G1341), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n684), .A2(G4), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n606), .B2(new_n684), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1348), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n824), .A2(G1341), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n821), .A2(new_n825), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n734), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n712), .A2(new_n831), .A3(new_n714), .A4(new_n732), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n735), .A2(new_n830), .A3(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n601), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n514), .B1(new_n837), .B2(KEYINPUT97), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(KEYINPUT97), .B2(new_n837), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n562), .A2(G93), .B1(G55), .B2(new_n523), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n547), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n606), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(new_n629), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n490), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n502), .A2(new_n504), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n498), .A2(KEYINPUT98), .A3(new_n499), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT98), .B1(new_n498), .B2(new_n499), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT99), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n500), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n857), .A4(new_n858), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n794), .A2(new_n795), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n786), .A2(KEYINPUT90), .A3(new_n787), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n788), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n754), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n800), .A2(KEYINPUT100), .A3(new_n753), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n872), .A2(new_n873), .A3(new_n766), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n766), .B1(new_n872), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n767), .ZN(new_n878));
  INV_X1    g453(.A(new_n866), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n873), .A3(new_n766), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n715), .A2(G142), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n479), .A2(G130), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n462), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n620), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(new_n720), .Z(new_n888));
  NAND3_X1  g463(.A1(new_n876), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n876), .A2(new_n881), .ZN(new_n892));
  INV_X1    g467(.A(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n890), .A3(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n856), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n856), .A2(new_n889), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n888), .B1(new_n876), .B2(new_n881), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n854), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n856), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n890), .B2(new_n889), .ZN(new_n904));
  INV_X1    g479(.A(new_n896), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT102), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n902), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G395));
  NAND2_X1  g486(.A1(new_n841), .A2(new_n590), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n844), .B(new_n613), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT103), .B1(new_n606), .B2(G299), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n567), .A2(new_n568), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n605), .A2(new_n915), .A3(new_n916), .A4(new_n563), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n606), .A2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n605), .A3(new_n563), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n913), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n913), .ZN(new_n926));
  INV_X1    g501(.A(new_n587), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n584), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT104), .B1(new_n927), .B2(new_n584), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n928), .A2(new_n929), .A3(new_n581), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n581), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n690), .A2(G303), .ZN(new_n933));
  OAI21_X1  g508(.A(G166), .B1(new_n687), .B2(new_n689), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n930), .A2(new_n934), .A3(new_n933), .A4(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT42), .Z(new_n939));
  XNOR2_X1  g514(.A(new_n926), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n912), .B1(new_n940), .B2(new_n590), .ZN(G295));
  OAI21_X1  g516(.A(new_n912), .B1(new_n940), .B2(new_n590), .ZN(G331));
  INV_X1    g517(.A(new_n843), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n549), .A2(new_n550), .B1(new_n839), .B2(new_n840), .ZN(new_n944));
  NOR2_X1   g519(.A1(G168), .A2(G171), .ZN(new_n945));
  AOI21_X1  g520(.A(G301), .B1(new_n532), .B2(new_n534), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(G301), .A2(new_n532), .A3(new_n534), .ZN(new_n948));
  NAND2_X1  g523(.A1(G168), .A2(G171), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n842), .A2(new_n843), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n921), .A3(new_n923), .ZN(new_n952));
  INV_X1    g527(.A(new_n925), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n936), .A2(KEYINPUT106), .A3(new_n937), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n938), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n956), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n955), .B2(new_n938), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n951), .A2(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n953), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n951), .A2(KEYINPUT41), .A3(new_n919), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n966), .A2(new_n961), .A3(new_n959), .A4(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n963), .A2(new_n968), .A3(KEYINPUT43), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n962), .B2(new_n963), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n963), .A2(new_n968), .A3(new_n971), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n974), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g550(.A1(new_n863), .A2(new_n857), .A3(new_n858), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n466), .A2(new_n469), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n473), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(G288), .A2(G1976), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT115), .Z(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  INV_X1    g560(.A(G1981), .ZN(new_n986));
  INV_X1    g561(.A(new_n579), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT114), .B(G86), .Z(new_n988));
  NAND2_X1  g563(.A1(new_n562), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n579), .A2(G1981), .A3(new_n580), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n581), .A2(new_n986), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n579), .B1(new_n562), .B2(new_n988), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n993), .B(KEYINPUT49), .C1(new_n986), .C2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n984), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n982), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n861), .A2(new_n865), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n494), .A2(G114), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(G2105), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n479), .A2(G126), .B1(new_n1005), .B2(new_n493), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n857), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n980), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1002), .B1(new_n1008), .B2(new_n999), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1001), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1971), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(KEYINPUT110), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1013));
  INV_X1    g588(.A(G2090), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n976), .A2(new_n1015), .A3(new_n980), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT110), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n998), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(KEYINPUT111), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G166), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1020), .A2(new_n1024), .A3(G8), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G288), .A2(new_n686), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(G1976), .A3(new_n688), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n982), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n995), .A2(new_n992), .A3(new_n982), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(G8), .A3(new_n981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT113), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(KEYINPUT113), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1037), .B(new_n1038), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n997), .B1(new_n1032), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1001), .A2(new_n743), .A3(new_n1009), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n976), .B2(new_n980), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1000), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n979), .B1(G164), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n743), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n979), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1015), .B1(new_n976), .B2(new_n980), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n1062), .A2(new_n1063), .A3(G2090), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1021), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1031), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1043), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1061), .A2(new_n1032), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1013), .A2(new_n808), .A3(new_n1016), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT116), .B(new_n1070), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(G168), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1025), .B1(KEYINPUT123), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(KEYINPUT123), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1073), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1075), .A2(new_n1074), .ZN(new_n1083));
  OAI211_X1 g658(.A(G8), .B(G286), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1080), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1069), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1079), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT62), .A3(new_n1084), .A4(new_n1081), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1044), .B1(new_n1068), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1032), .A2(new_n1067), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(G168), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1020), .A2(G8), .A3(new_n1024), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1031), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1020), .A2(new_n1101), .A3(new_n1024), .A4(G8), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1043), .A2(new_n1095), .A3(new_n1093), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1001), .A2(new_n1009), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n816), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT57), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT57), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n915), .A2(new_n563), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(G299), .A2(new_n1110), .A3(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n981), .A2(KEYINPUT119), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n976), .A2(new_n979), .A3(new_n1118), .A4(new_n980), .ZN(new_n1119));
  AOI21_X1  g694(.A(G2067), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1048), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1120), .A2(KEYINPUT120), .B1(new_n1121), .B2(G1348), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1107), .A2(new_n1108), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n606), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1116), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT58), .B(G1341), .Z(new_n1129));
  NAND3_X1  g704(.A1(new_n1117), .A2(new_n1119), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1001), .A2(new_n1131), .A3(new_n1009), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n552), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1133), .B2(new_n552), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1128), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1137), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(KEYINPUT59), .A3(new_n1135), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1116), .A2(new_n1125), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND4_X1   g719(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n606), .A2(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n606), .A2(KEYINPUT122), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1122), .A2(new_n1123), .A3(new_n1149), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1148), .B(new_n1150), .C1(new_n1151), .C2(new_n1146), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1127), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1032), .A2(new_n1067), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1002), .A2(new_n1046), .A3(G2078), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n861), .A2(new_n980), .A3(new_n865), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(KEYINPUT107), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n999), .B1(new_n1157), .B2(KEYINPUT107), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1001), .B(new_n1156), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(G301), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1059), .A2(new_n1060), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1155), .A2(G301), .A3(new_n1055), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT54), .B(new_n1165), .C1(new_n1166), .C2(G301), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1089), .A2(new_n1084), .A3(new_n1081), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1154), .A2(new_n1164), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1092), .B(new_n1105), .C1(new_n1153), .C2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1158), .A2(new_n1159), .A3(new_n1002), .ZN(new_n1171));
  INV_X1    g746(.A(G1986), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n588), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n588), .A2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n753), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n1131), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n766), .B(G2067), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1171), .A2(KEYINPUT109), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT109), .B1(new_n1171), .B2(new_n1179), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1171), .A2(new_n1131), .A3(new_n754), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT108), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n720), .B(new_n726), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1185), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1176), .A2(new_n1182), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1170), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .A4(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1171), .B1(new_n753), .B2(new_n1179), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT126), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1171), .B(new_n1194), .C1(new_n753), .C2(new_n1179), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT47), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1171), .A2(new_n1131), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT46), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1191), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1171), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n721), .A2(new_n726), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT125), .Z(new_n1205));
  NAND3_X1  g780(.A1(new_n1182), .A2(new_n1184), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n767), .A2(new_n769), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1203), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1188), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(G319), .ZN(new_n1212));
  OR2_X1    g786(.A1(G227), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g787(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n1214), .A2(new_n647), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G229), .A2(new_n1216), .ZN(new_n1217));
  NOR3_X1   g791(.A1(new_n897), .A2(new_n854), .A3(new_n901), .ZN(new_n1218));
  AOI21_X1  g792(.A(KEYINPUT102), .B1(new_n906), .B2(new_n907), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g794(.A1(new_n1220), .A2(new_n974), .ZN(G308));
  OAI221_X1 g795(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .C1(new_n972), .C2(new_n973), .ZN(G225));
endmodule


