//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(new_n460), .A3(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OR3_X1    g045(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(KEYINPUT3), .B(G2104), .Z(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(G2105), .B1(G101), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n482), .A2(G100), .A3(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n465), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(G100), .B2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(G2104), .A3(new_n485), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n469), .A2(new_n481), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n466), .A2(new_n468), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(G2105), .A3(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n487), .B1(new_n490), .B2(G124), .ZN(G162));
  NAND4_X1  g066(.A1(new_n488), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n493), .A2(new_n465), .A3(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n465), .B2(G114), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n494), .A2(G2104), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT72), .B1(new_n474), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT3), .B(G2104), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n469), .B2(new_n499), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n488), .A2(G138), .A3(new_n465), .A4(new_n464), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT4), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n498), .B1(new_n508), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n518), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n525), .A2(G88), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n519), .ZN(new_n531));
  OAI211_X1 g106(.A(G543), .B(new_n531), .C1(new_n526), .C2(new_n513), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n530), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NOR2_X1   g111(.A1(new_n516), .A2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT6), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n539), .A2(G51), .A3(G543), .A4(new_n531), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n521), .A2(new_n523), .A3(G63), .A4(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT7), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT5), .B(G543), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n539), .A2(G89), .A3(new_n531), .A4(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n540), .A2(new_n546), .A3(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n524), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n526), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n539), .A2(G90), .A3(new_n531), .A4(new_n547), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n539), .A2(G52), .A3(G543), .A4(new_n531), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G171));
  NOR2_X1   g132(.A1(new_n518), .A2(new_n519), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT74), .B(G81), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(new_n547), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n524), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(new_n526), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n539), .A2(G43), .A3(G543), .A4(new_n531), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G188));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n558), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n532), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n539), .A2(G91), .A3(new_n531), .A4(new_n547), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n547), .A2(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(G299));
  NAND2_X1  g161(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  OAI21_X1  g166(.A(G651), .B1(new_n547), .B2(G74), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT78), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n533), .A2(G49), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n525), .A2(G87), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n524), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n525), .A2(G86), .B1(new_n526), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n533), .A2(G48), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n547), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(new_n526), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n539), .A2(G47), .A3(G543), .A4(new_n531), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n539), .A2(G85), .A3(new_n531), .A4(new_n547), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(KEYINPUT80), .B(new_n605), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G54), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n547), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OAI22_X1  g193(.A1(new_n532), .A2(new_n617), .B1(new_n618), .B2(new_n514), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n531), .B(new_n547), .C1(new_n526), .C2(new_n513), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(G868), .B2(new_n625), .ZN(G284));
  OAI21_X1  g201(.A(new_n616), .B1(G868), .B2(new_n625), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n585), .A2(new_n580), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n578), .B2(new_n576), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n625), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n490), .A2(G123), .ZN(new_n639));
  INV_X1    g214(.A(new_n469), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G135), .ZN(new_n641));
  OR2_X1    g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(G2096), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n503), .A2(new_n477), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XOR2_X1   g226(.A(KEYINPUT13), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n679), .A2(KEYINPUT17), .A3(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n676), .B1(new_n679), .B2(KEYINPUT17), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n680), .A2(new_n681), .A3(new_n675), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n692), .B1(new_n687), .B2(new_n690), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1991), .ZN(new_n698));
  INV_X1    g273(.A(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1971), .Z(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT87), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n709), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G24), .B(G290), .S(G16), .Z(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1986), .Z(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  INV_X1    g300(.A(G131), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT85), .B1(new_n469), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G119), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n465), .A2(G107), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n727), .B1(new_n728), .B2(new_n489), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n726), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(new_n724), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n721), .A2(new_n723), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT88), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n720), .B2(new_n718), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT36), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(G29), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT97), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n724), .A2(G26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n490), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n640), .A2(G140), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(new_n724), .ZN(new_n756));
  MUX2_X1   g331(.A(new_n749), .B(new_n756), .S(KEYINPUT28), .Z(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n724), .A2(G33), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n465), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT89), .Z(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n477), .A2(G103), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  INV_X1    g341(.A(G139), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n469), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n760), .B1(new_n770), .B2(new_n724), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G2072), .Z(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n724), .B1(new_n773), .B2(G28), .ZN(new_n775));
  AND2_X1   g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NOR2_X1   g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G168), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G16), .B2(G21), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(new_n724), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n479), .B2(new_n724), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2084), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n625), .B2(G16), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1348), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1348), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n567), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n644), .A2(new_n724), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n796), .B(new_n798), .C1(new_n781), .C2(new_n780), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n783), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n747), .A2(new_n748), .A3(new_n759), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n710), .A2(G5), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G171), .B2(new_n710), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1961), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n710), .A2(G20), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n806), .B(new_n807), .C1(G299), .C2(G16), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n724), .A2(G27), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n724), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2078), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n801), .A2(new_n805), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n640), .A2(G141), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT91), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n490), .A2(G129), .ZN(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT26), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n821), .A2(new_n822), .B1(G105), .B2(new_n477), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT92), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n724), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT93), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G29), .B2(G32), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT27), .Z(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(G1996), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(G1996), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n740), .B(new_n814), .C1(new_n830), .C2(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  XNOR2_X1  g408(.A(KEYINPUT98), .B(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n625), .A2(G559), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n539), .A2(G93), .A3(new_n531), .A4(new_n547), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n547), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n838), .B1(new_n532), .B2(new_n839), .C1(new_n604), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n566), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n834), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n834), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n479), .B(new_n644), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(G162), .Z(new_n849));
  XNOR2_X1  g424(.A(G164), .B(new_n755), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n769), .B1(new_n825), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n825), .B2(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  INV_X1    g428(.A(new_n850), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n770), .B1(new_n854), .B2(new_n824), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n824), .B2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n853), .B2(new_n852), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n490), .A2(G130), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n640), .A2(G142), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n465), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n733), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n651), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n651), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n858), .A2(new_n869), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n849), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  INV_X1    g449(.A(new_n849), .ZN(new_n875));
  INV_X1    g450(.A(new_n867), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n870), .B(new_n875), .C1(new_n876), .C2(new_n858), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(G395));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n624), .A2(new_n623), .ZN(new_n882));
  INV_X1    g457(.A(new_n619), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n630), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(G299), .A2(new_n625), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n630), .A2(new_n884), .ZN(new_n890));
  NOR2_X1   g465(.A1(G299), .A2(new_n625), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n889), .B1(new_n894), .B2(new_n881), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n842), .B(new_n635), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n895), .A2(KEYINPUT103), .A3(new_n896), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n901), .B(new_n903), .Z(new_n904));
  XNOR2_X1  g479(.A(G303), .B(G305), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n613), .A2(new_n614), .A3(G288), .ZN(new_n907));
  AOI21_X1  g482(.A(G288), .B1(new_n613), .B2(new_n614), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G290), .A2(new_n706), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n613), .A2(new_n614), .A3(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n902), .B2(KEYINPUT42), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n904), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(new_n914), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n915), .A2(new_n916), .A3(G868), .A4(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(G868), .A3(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(G868), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT105), .B1(new_n841), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(G295));
  OAI21_X1  g497(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(G331));
  NOR2_X1   g498(.A1(G168), .A2(new_n556), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(G301), .B2(G168), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(new_n842), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n842), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n887), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n925), .A2(new_n929), .A3(new_n842), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n925), .B2(new_n842), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n925), .A2(new_n842), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n913), .B(new_n928), .C1(new_n895), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n934), .B2(KEYINPUT108), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n930), .A2(new_n931), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(new_n885), .B2(new_n886), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n881), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n936), .A2(new_n926), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n913), .A4(new_n928), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n935), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(new_n928), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n913), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(new_n928), .C1(new_n895), .C2(new_n933), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n935), .A3(new_n947), .A4(new_n944), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT109), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n936), .A2(new_n887), .A3(new_n926), .ZN(new_n958));
  INV_X1    g533(.A(new_n894), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n926), .A2(new_n927), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n950), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n935), .A2(new_n944), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n963), .B2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT110), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n954), .A2(new_n956), .A3(new_n964), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n945), .A2(new_n953), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(KEYINPUT43), .B2(new_n963), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n957), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(new_n973), .A3(KEYINPUT111), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(G164), .B2(G1384), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT112), .B(G40), .ZN(new_n981));
  AND4_X1   g556(.A1(new_n471), .A2(new_n472), .A3(new_n478), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n733), .A2(new_n735), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n733), .A2(new_n735), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n699), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n825), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n754), .B(G2067), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n984), .A2(KEYINPUT113), .A3(G1996), .A4(new_n824), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n984), .A2(new_n824), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(new_n699), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(G290), .B(G1986), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n988), .B(new_n997), .C1(new_n984), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT4), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n510), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n506), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n1000), .C1(new_n1003), .C2(new_n498), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n980), .A2(new_n1004), .A3(new_n982), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n781), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n1007));
  INV_X1    g582(.A(new_n506), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n511), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n498), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n982), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1006), .B1(G2084), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G8), .A3(G286), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n1017), .B(KEYINPUT121), .Z(new_n1018));
  OAI211_X1 g593(.A(new_n1006), .B(G168), .C1(G2084), .C2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT122), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1019), .A2(new_n1024), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n982), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1030));
  NOR3_X1   g605(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G1961), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1005), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2078), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n980), .A2(new_n1004), .A3(KEYINPUT114), .A4(new_n982), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n980), .A2(new_n1004), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(G2078), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(G40), .A3(G160), .A4(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1029), .B(new_n556), .C1(new_n1040), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1033), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1043), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT124), .B1(new_n1047), .B2(G171), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n982), .A3(new_n1042), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1040), .A2(G301), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1040), .A2(new_n1053), .A3(G301), .A4(new_n1050), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT125), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  AND4_X1   g632(.A1(G301), .A2(new_n1045), .A3(new_n1046), .A4(new_n1043), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1040), .B2(new_n1050), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1015), .A2(G2090), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G303), .A2(G8), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n1067), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1011), .A2(new_n982), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n706), .A2(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(G8), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G305), .A2(G1981), .ZN(new_n1076));
  INV_X1    g651(.A(G1981), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n600), .B2(new_n601), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT115), .B(new_n1081), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1069), .A3(G8), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1072), .A2(new_n1075), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT116), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1072), .A2(new_n1086), .A3(new_n1083), .A4(new_n1075), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1066), .A2(new_n1068), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1060), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1092));
  XNOR2_X1  g667(.A(G299), .B(KEYINPUT57), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n980), .A2(new_n1004), .A3(new_n982), .A4(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1069), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1015), .A2(new_n1098), .B1(new_n1099), .B2(new_n758), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(new_n884), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1093), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1094), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1097), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT119), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n980), .A2(new_n1004), .A3(new_n699), .A4(new_n982), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1069), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1115), .B2(new_n567), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1111), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n566), .B(new_n1117), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1107), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1015), .A2(new_n1098), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1099), .A2(new_n758), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n884), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n1122), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n625), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1100), .A2(new_n1127), .A3(KEYINPUT60), .A4(new_n884), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1100), .A2(KEYINPUT60), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1104), .B1(new_n1120), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1090), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1047), .A2(G171), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1029), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1047), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(KEYINPUT54), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1056), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1059), .A2(new_n1066), .A3(new_n1068), .A4(new_n1088), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1027), .B2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1028), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1083), .A2(new_n1073), .A3(new_n706), .ZN(new_n1146));
  OAI211_X1 g721(.A(G8), .B(new_n1069), .C1(new_n1146), .C2(new_n1076), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1068), .B2(new_n1084), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1143), .B2(KEYINPUT62), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1016), .A2(G8), .A3(G168), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1066), .A2(new_n1068), .A3(new_n1088), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n1151), .B2(KEYINPUT117), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(KEYINPUT117), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1067), .A2(KEYINPUT118), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1063), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1063), .A2(new_n1154), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1084), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1155), .A2(new_n1150), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1149), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n999), .B1(new_n1145), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n985), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n997), .A2(new_n1165), .A3(new_n988), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n989), .B(KEYINPUT46), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n984), .B1(new_n991), .B2(new_n824), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(KEYINPUT126), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(KEYINPUT126), .B2(new_n1168), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT47), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n997), .A2(new_n986), .B1(G2067), .B2(new_n754), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1166), .B(new_n1171), .C1(new_n984), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1162), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(G319), .ZN(new_n1176));
  INV_X1    g750(.A(new_n670), .ZN(new_n1177));
  NOR4_X1   g751(.A1(G229), .A2(new_n1176), .A3(new_n1177), .A4(G227), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1178), .A2(new_n878), .A3(new_n972), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


