//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n202), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n210), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(new_n211), .B1(G20), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(G20), .B1(G33), .B2(G283), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G97), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT87), .ZN(new_n252));
  AND3_X1   g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n249), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(KEYINPUT20), .B(new_n248), .C1(new_n253), .C2(new_n254), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n257), .A2(new_n258), .B1(new_n247), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT69), .B1(new_n246), .B2(new_n211), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT76), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n269), .B2(new_n263), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n259), .A2(G33), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n268), .A2(new_n271), .A3(G116), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G303), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n283), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n277), .A2(KEYINPUT82), .A3(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT82), .B1(new_n277), .B2(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n276), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n280), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT5), .B(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  INV_X1    g0097(.A(new_n211), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n294), .A2(G270), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n275), .B1(new_n290), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n274), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT21), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n290), .A2(G179), .A3(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n274), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n274), .A2(KEYINPUT21), .A3(new_n302), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n305), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n290), .A2(new_n301), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G200), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n290), .B2(new_n301), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n313), .A2(new_n274), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT3), .B(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n283), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G222), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n319), .A2(new_n320), .B1(new_n321), .B2(new_n318), .ZN(new_n322));
  INV_X1    g0122(.A(G223), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n279), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n289), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G41), .ZN(new_n327));
  AOI21_X1  g0127(.A(G1), .B1(new_n327), .B2(new_n291), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n300), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n289), .A2(new_n328), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(G226), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n314), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT79), .Z(new_n335));
  NOR2_X1   g0135(.A1(new_n269), .A2(new_n263), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n203), .A2(G20), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT71), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT70), .A2(G58), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT8), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n250), .A2(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G20), .A2(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n336), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G50), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n259), .B2(G20), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n266), .A2(new_n349), .B1(new_n348), .B2(new_n261), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(KEYINPUT9), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT78), .B1(new_n333), .B2(G190), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n335), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT10), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT10), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n335), .A2(new_n359), .A3(new_n351), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT73), .B1(new_n333), .B2(G169), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT72), .B(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n333), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n352), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT8), .B(G58), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n345), .B1(new_n212), .B2(new_n321), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n341), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n372), .B(new_n373), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n336), .B1(new_n321), .B2(new_n261), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n259), .A2(G20), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n268), .A2(new_n271), .A3(G77), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(KEYINPUT77), .A3(new_n382), .ZN(new_n386));
  OR2_X1    g0186(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n318), .B1(new_n219), .B2(new_n324), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n289), .C1(G107), .C2(new_n318), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n330), .B1(G244), .B2(new_n331), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(G190), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n385), .A2(new_n386), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n363), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n275), .B2(new_n395), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n383), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n361), .A2(new_n369), .A3(new_n397), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n283), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT80), .B(new_n403), .C1(new_n404), .C2(new_n279), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT80), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n387), .A2(G226), .A3(new_n388), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G232), .A2(G1698), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n279), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n403), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n411), .A3(new_n289), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n330), .B1(G238), .B2(new_n331), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT81), .B1(new_n418), .B2(new_n312), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n412), .A2(new_n416), .A3(new_n413), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n412), .B2(new_n413), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT81), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(G190), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n264), .A2(new_n265), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n341), .A2(G77), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n344), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT11), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n261), .A2(new_n218), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT12), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(KEYINPUT11), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND4_X1   g0234(.A1(G68), .A2(new_n268), .A3(new_n271), .A4(new_n381), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n422), .B2(new_n314), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n434), .A2(new_n435), .ZN(new_n440));
  OAI21_X1  g0240(.A(G169), .B1(new_n420), .B2(new_n421), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n441), .A2(KEYINPUT14), .B1(new_n418), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n418), .B2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n340), .A2(new_n381), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n270), .A2(new_n448), .B1(new_n260), .B2(new_n340), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI221_X1 g0251(.A(KEYINPUT85), .B1(new_n260), .B2(new_n340), .C1(new_n270), .C2(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G58), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n218), .ZN(new_n455));
  OAI21_X1  g0255(.A(G20), .B1(new_n455), .B2(new_n202), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n344), .A2(G159), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n277), .A2(KEYINPUT82), .A3(G33), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(G20), .B1(new_n462), .B2(new_n276), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT7), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n218), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n277), .A2(G33), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT7), .B1(new_n467), .B2(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n458), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n426), .B1(new_n469), .B2(KEYINPUT16), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT16), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  AOI21_X1  g0272(.A(G20), .B1(new_n276), .B2(new_n278), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(KEYINPUT7), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT83), .B(new_n464), .C1(new_n318), .C2(G20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n250), .A2(KEYINPUT84), .A3(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n278), .A2(KEYINPUT84), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n276), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n464), .A2(G20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n218), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n471), .B1(new_n482), .B2(new_n458), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n453), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n283), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n485), .A2(new_n287), .B1(new_n250), .B2(new_n220), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n289), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n331), .A2(G232), .B1(new_n300), .B2(new_n328), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n275), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G226), .A2(G1698), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n389), .B2(new_n323), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(new_n467), .B1(G33), .B2(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n298), .A2(new_n299), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n398), .B(new_n488), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n484), .A2(KEYINPUT18), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT18), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n451), .A2(new_n452), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n212), .B1(new_n466), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT83), .B1(new_n501), .B2(new_n464), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n473), .A2(new_n472), .A3(KEYINPUT7), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n481), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G68), .ZN(new_n505));
  INV_X1    g0305(.A(new_n458), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT16), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n287), .A2(new_n464), .A3(new_n212), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n468), .A3(G68), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT16), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n336), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n499), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n488), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n486), .B2(new_n289), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n494), .B1(new_n514), .B2(new_n275), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n498), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n458), .B1(new_n504), .B2(G68), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n336), .B(new_n510), .C1(new_n518), .C2(KEYINPUT16), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n487), .A2(new_n312), .A3(new_n488), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n514), .B2(G200), .ZN(new_n521));
  AND4_X1   g0321(.A1(KEYINPUT17), .A2(new_n519), .A3(new_n499), .A4(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT17), .B1(new_n484), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n402), .A2(new_n447), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n212), .B2(G107), .ZN(new_n530));
  INV_X1    g0330(.A(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n250), .A2(new_n247), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n535), .B2(G20), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n220), .A2(G20), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT22), .B1(new_n318), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n220), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n467), .A2(new_n212), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n528), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n318), .A2(new_n537), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n530), .A2(new_n532), .B1(new_n534), .B2(new_n212), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n542), .A2(new_n545), .A3(new_n546), .A4(new_n528), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n336), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT89), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT89), .B(new_n336), .C1(new_n543), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n260), .A2(KEYINPUT91), .A3(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT90), .B(KEYINPUT25), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT91), .B1(new_n260), .B2(G107), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(KEYINPUT91), .C1(G107), .C2(new_n260), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n260), .B(new_n272), .C1(new_n269), .C2(new_n263), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n531), .C2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G257), .A2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n389), .B2(new_n221), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n467), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n493), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n294), .A2(G264), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n296), .A2(new_n300), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n442), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n294), .A2(G264), .B1(new_n296), .B2(new_n300), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n564), .A2(new_n467), .B1(G33), .B2(G294), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n493), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n275), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n567), .B2(new_n570), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n573), .B(G190), .C1(new_n574), .C2(new_n493), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(new_n561), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n562), .A2(new_n578), .B1(new_n552), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n261), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n559), .B2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n531), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n583), .A2(new_n531), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n589), .B2(KEYINPUT6), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n344), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n474), .A2(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n531), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n585), .B1(new_n593), .B2(new_n336), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n318), .A2(G250), .A3(G1698), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G283), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT4), .A2(G244), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n596), .C1(new_n319), .C2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n387), .A2(G244), .A3(new_n388), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT4), .B1(new_n467), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n289), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n294), .A2(G257), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n569), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(new_n314), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(G190), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n594), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n275), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n601), .A2(new_n569), .A3(new_n363), .A4(new_n602), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n593), .A2(new_n336), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n585), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n377), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  INV_X1    g0413(.A(new_n559), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT86), .B1(new_n377), .B2(new_n559), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n467), .A2(new_n212), .A3(G68), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n341), .A2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n212), .B1(new_n403), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n588), .A2(new_n220), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n426), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n260), .B1(new_n375), .B2(new_n376), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n300), .A2(new_n292), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n292), .A2(new_n221), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n493), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n387), .A2(G238), .A3(new_n388), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G244), .A2(G1698), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n534), .B1(new_n634), .B2(new_n467), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n631), .B1(new_n635), .B2(new_n493), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G169), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n631), .B(new_n398), .C1(new_n635), .C2(new_n493), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n628), .A2(new_n630), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n283), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n535), .B1(new_n642), .B2(new_n287), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n289), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G190), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n559), .A2(new_n220), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n624), .A2(new_n646), .A3(new_n625), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n636), .A2(G200), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n317), .A2(new_n526), .A3(new_n582), .A4(new_n651), .ZN(G372));
  NAND3_X1  g0452(.A1(new_n439), .A2(new_n383), .A3(new_n400), .ZN(new_n653));
  AOI211_X1 g0453(.A(new_n523), .B(new_n522), .C1(new_n653), .C2(new_n446), .ZN(new_n654));
  INV_X1    g0454(.A(new_n517), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n361), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n369), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n603), .A2(new_n275), .ZN(new_n658));
  INV_X1    g0458(.A(new_n608), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n594), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n638), .B(KEYINPUT92), .C1(new_n644), .C2(new_n275), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT92), .B1(new_n637), .B2(new_n638), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n627), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(new_n646), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n626), .A2(KEYINPUT93), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT93), .B1(new_n626), .B2(new_n666), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n648), .B(new_n645), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n660), .A2(new_n664), .A3(new_n665), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n650), .B2(new_n610), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n670), .A2(new_n671), .A3(new_n664), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n552), .A2(new_n581), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n673), .A2(new_n610), .A3(new_n606), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n309), .A2(new_n308), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n560), .B1(new_n550), .B2(new_n551), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n675), .B(new_n305), .C1(new_n676), .C2(new_n577), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n664), .A2(new_n669), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n526), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT94), .Z(G369));
  NAND3_X1  g0484(.A1(new_n259), .A2(new_n212), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n274), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n317), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n310), .A2(new_n274), .A3(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT95), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT95), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n696), .A3(new_n693), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(G330), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n690), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n582), .B1(new_n676), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n577), .B1(new_n552), .B2(new_n561), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n310), .A2(new_n700), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n582), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n700), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT96), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(KEYINPUT96), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n705), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n208), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n622), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n216), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n571), .A2(new_n644), .A3(new_n601), .A4(new_n602), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n306), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n575), .A2(new_n636), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n601), .A2(new_n602), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n307), .A3(KEYINPUT30), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n571), .A2(new_n398), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n311), .A3(new_n636), .A4(new_n603), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n690), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n651), .A2(new_n582), .A3(new_n317), .A4(new_n700), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n723), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n664), .B(KEYINPUT97), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT26), .B1(new_n678), .B2(new_n610), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n660), .A2(new_n665), .A3(new_n640), .A4(new_n649), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n702), .A2(new_n310), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n673), .A2(new_n610), .A3(new_n606), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n742), .A2(new_n743), .A3(new_n678), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n700), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT98), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(KEYINPUT98), .B(new_n700), .C1(new_n741), .C2(new_n744), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n690), .B1(new_n672), .B2(new_n680), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT29), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n737), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n722), .B1(new_n753), .B2(G1), .ZN(G364));
  AND2_X1   g0554(.A1(new_n695), .A2(new_n697), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n212), .A2(G13), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n259), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n717), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n756), .A2(new_n699), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT99), .Z(new_n762));
  NOR2_X1   g0562(.A1(new_n716), .A2(new_n279), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G355), .A2(new_n763), .B1(new_n247), .B2(new_n716), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n244), .A2(new_n291), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n467), .A2(new_n716), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n216), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n211), .B1(G20), .B2(new_n275), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n717), .B(new_n759), .C1(new_n768), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n212), .A2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n314), .A2(G179), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G283), .A2(new_n779), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n783), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n212), .A2(new_n312), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n777), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n279), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT100), .Z(new_n793));
  NAND3_X1  g0593(.A1(new_n398), .A2(new_n314), .A3(new_n789), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n788), .B(new_n793), .C1(G322), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n398), .A2(G20), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  INV_X1    g0601(.A(new_n776), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n363), .A2(new_n802), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n797), .A2(new_n312), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G326), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n806), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n808), .A2(new_n348), .B1(new_n321), .B2(new_n804), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G58), .B2(new_n795), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n318), .B1(new_n778), .B2(new_n531), .C1(new_n220), .C2(new_n790), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n781), .B2(new_n812), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n583), .C2(new_n787), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n811), .B(new_n815), .C1(G68), .C2(new_n798), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n796), .A2(new_n807), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n771), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n774), .B1(new_n775), .B2(new_n817), .C1(new_n755), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n762), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(G396));
  NOR2_X1   g0622(.A1(new_n401), .A2(new_n690), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n383), .A2(new_n690), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n397), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n401), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n751), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n670), .A2(new_n671), .A3(new_n664), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n700), .C1(new_n744), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n737), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n760), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n737), .A3(new_n829), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n795), .A2(G143), .B1(G159), .B2(new_n803), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n808), .B2(new_n836), .C1(new_n343), .C2(new_n799), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n779), .A2(G68), .ZN(new_n839));
  INV_X1    g0639(.A(new_n790), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G50), .A2(new_n840), .B1(new_n782), .B2(G132), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n287), .B1(G58), .B2(new_n786), .ZN(new_n842));
  AND4_X1   g0642(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n798), .A2(G283), .B1(G116), .B2(new_n803), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n784), .B2(new_n794), .C1(new_n791), .C2(new_n808), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n787), .A2(new_n583), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n279), .B1(new_n781), .B2(new_n801), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n779), .A2(G87), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n531), .B2(new_n790), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n772), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n775), .A2(new_n770), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n760), .C1(G77), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n826), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n769), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n834), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  AOI211_X1 g0658(.A(new_n247), .B(new_n214), .C1(new_n590), .C2(KEYINPUT35), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n590), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OR3_X1    g0661(.A1(new_n216), .A2(new_n321), .A3(new_n455), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n201), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n259), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n509), .B2(new_n506), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n499), .B1(new_n511), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n688), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n517), .B2(new_n524), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n512), .A2(new_n515), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n512), .A2(new_n868), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n519), .A2(new_n499), .A3(new_n521), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n867), .A2(new_n515), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n880), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n871), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n871), .C1(new_n878), .C2(new_n885), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n880), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT104), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n519), .A2(new_n499), .A3(new_n521), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n496), .B1(new_n519), .B2(new_n499), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n897), .A2(new_n877), .A3(new_n874), .A4(new_n873), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n887), .B(new_n870), .C1(new_n894), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n873), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n873), .B1(new_n517), .B2(new_n524), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n891), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n418), .A2(new_n444), .A3(G169), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n911), .B(new_n912), .C1(new_n442), .C2(new_n418), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n440), .A3(new_n700), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n890), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n655), .A2(new_n688), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n888), .A2(new_n889), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT103), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n823), .B1(new_n751), .B2(new_n826), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n437), .B1(new_n424), .B2(new_n419), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n440), .B(new_n690), .C1(new_n921), .C2(new_n913), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n440), .A2(new_n690), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n439), .A2(new_n446), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n919), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n823), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n829), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT103), .A3(new_n925), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n918), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n916), .A2(new_n917), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n750), .A2(new_n526), .A3(new_n752), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n657), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n932), .B(new_n934), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n735), .A2(new_n736), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n925), .A2(new_n936), .A3(new_n826), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n894), .A2(new_n900), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n938), .B2(new_n871), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n939), .B2(new_n901), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n898), .A2(new_n899), .B1(new_n902), .B2(KEYINPUT37), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n887), .B1(new_n943), .B2(new_n907), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n889), .A2(new_n944), .ZN(new_n945));
  AND4_X1   g0745(.A1(KEYINPUT40), .A2(new_n925), .A3(new_n936), .A4(new_n826), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n526), .A2(new_n936), .ZN(new_n949));
  OAI21_X1  g0749(.A(G330), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n935), .A2(new_n951), .B1(new_n259), .B2(new_n757), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n935), .A2(new_n951), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n865), .B1(new_n952), .B2(new_n953), .ZN(G367));
  INV_X1    g0754(.A(new_n766), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n773), .B1(new_n208), .B2(new_n377), .C1(new_n233), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n760), .ZN(new_n957));
  INV_X1    g0757(.A(new_n201), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n795), .A2(G150), .B1(new_n958), .B2(new_n803), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n808), .B2(new_n960), .C1(new_n812), .C2(new_n799), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n787), .A2(new_n218), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n318), .B1(new_n781), .B2(new_n836), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n790), .A2(new_n454), .B1(new_n778), .B2(new_n321), .ZN(new_n964));
  NOR4_X1   g0764(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n806), .A2(G311), .B1(new_n795), .B2(G303), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n784), .B2(new_n799), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n840), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n790), .B2(new_n247), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(new_n531), .C2(new_n787), .ZN(new_n971));
  INV_X1    g0771(.A(G283), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n804), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n779), .A2(G97), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n782), .A2(G317), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n975), .A3(new_n287), .ZN(new_n976));
  NOR4_X1   g0776(.A1(new_n967), .A2(new_n971), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n965), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  AOI21_X1  g0779(.A(new_n957), .B1(new_n979), .B2(new_n772), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n667), .A2(new_n668), .A3(new_n700), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n679), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n664), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n771), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n708), .B1(new_n704), .B2(new_n707), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT109), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n698), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(new_n753), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n606), .B(new_n610), .C1(new_n594), .C2(new_n700), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n660), .A2(new_n690), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n714), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT45), .B1(new_n714), .B2(new_n994), .ZN(new_n998));
  INV_X1    g0798(.A(new_n994), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n712), .A2(new_n713), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n997), .A2(new_n998), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n699), .A3(new_n704), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n705), .B1(new_n1002), .B2(new_n1003), .C1(new_n997), .C2(new_n998), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n991), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n753), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n717), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n759), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n999), .B2(new_n708), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT42), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n582), .A4(new_n707), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT107), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n610), .B1(new_n992), .B2(new_n703), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n700), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n982), .A2(new_n983), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT108), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1021), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1030), .A2(new_n1031), .B1(new_n705), .B2(new_n999), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1031), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n705), .A2(new_n999), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n1029), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n985), .B1(new_n1011), .B2(new_n1036), .ZN(G387));
  OR2_X1    g0837(.A1(new_n704), .A2(new_n818), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n763), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1039), .A2(new_n719), .B1(G107), .B2(new_n208), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n237), .A2(new_n291), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n719), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n370), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n955), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n773), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n760), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G159), .A2(new_n806), .B1(new_n798), .B2(new_n340), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n612), .A2(new_n786), .B1(G68), .B2(new_n803), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n840), .A2(G77), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n974), .C1(new_n343), .C2(new_n781), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n287), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n795), .A2(G50), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G116), .A2(new_n779), .B1(new_n782), .B2(G326), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n787), .A2(new_n972), .B1(new_n790), .B2(new_n784), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n795), .A2(G317), .B1(G303), .B2(new_n803), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT111), .B(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n808), .B2(new_n1061), .C1(new_n801), .C2(new_n799), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n287), .B(new_n1058), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1057), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n775), .B1(new_n1069), .B2(KEYINPUT112), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1050), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n990), .A2(new_n759), .B1(new_n1038), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n990), .A2(new_n753), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n717), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n990), .A2(new_n753), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  AND2_X1   g0877(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n999), .A2(new_n771), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n773), .B1(new_n583), .B2(new_n208), .C1(new_n241), .C2(new_n955), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n760), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n806), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n798), .A2(G303), .B1(G116), .B2(new_n786), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n790), .A2(new_n972), .B1(new_n781), .B2(new_n1061), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n318), .B(new_n1088), .C1(G107), .C2(new_n779), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n784), .B2(new_n804), .C1(new_n1085), .C2(KEYINPUT114), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n806), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n799), .A2(new_n201), .B1(new_n370), .B2(new_n804), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n848), .B1(new_n218), .B2(new_n790), .C1(new_n960), .C2(new_n781), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n786), .A2(G77), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n467), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1087), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1081), .B1(new_n1098), .B2(new_n772), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1078), .A2(new_n759), .B1(new_n1079), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1074), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1007), .A2(new_n1102), .A3(new_n717), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(KEYINPUT115), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT115), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n718), .B1(new_n1078), .B2(new_n991), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n1102), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1104), .B2(new_n1107), .ZN(G390));
  NAND3_X1  g0908(.A1(new_n737), .A2(new_n826), .A3(new_n925), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n747), .A2(new_n748), .A3(new_n928), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n825), .A2(new_n401), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n925), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n915), .B1(new_n889), .B2(new_n944), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n915), .B1(new_n929), .B2(new_n925), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n890), .B2(new_n910), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1110), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n1109), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n526), .A2(new_n737), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n933), .A2(new_n657), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n737), .A2(new_n826), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n926), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n920), .B1(new_n1126), .B2(new_n1109), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(new_n1109), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT116), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1122), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1118), .B(new_n1121), .C1(new_n1131), .C2(KEYINPUT116), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n717), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1122), .B2(new_n758), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1118), .A2(new_n1121), .A3(KEYINPUT117), .A4(new_n759), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n760), .B1(new_n340), .B2(new_n852), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n806), .A2(G283), .B1(G97), .B2(new_n803), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n531), .B2(new_n799), .C1(new_n247), .C2(new_n794), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n318), .B1(new_n840), .B2(G87), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n782), .A2(G294), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n839), .A3(new_n1095), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n318), .B1(new_n781), .B2(new_n1147), .C1(new_n201), .C2(new_n778), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n806), .B2(G128), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n840), .A2(G150), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1150), .A2(KEYINPUT53), .B1(G159), .B2(new_n786), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(KEYINPUT53), .C2(new_n1150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n795), .A2(G132), .B1(new_n803), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n836), .B2(new_n799), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1143), .A2(new_n1146), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1141), .B1(new_n1157), .B2(new_n772), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n890), .A2(new_n910), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n770), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1136), .A2(new_n1140), .A3(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n723), .B1(new_n945), .B2(new_n946), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n352), .A2(new_n868), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n361), .B2(new_n369), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1164), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1167), .B(new_n368), .C1(new_n358), .C2(new_n360), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1170), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n942), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n942), .B2(new_n1163), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n932), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT40), .B1(new_n918), .B2(new_n937), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n947), .A2(G330), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n942), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n929), .A2(new_n925), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(new_n919), .B1(new_n888), .B2(new_n889), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1184), .A2(new_n930), .B1(new_n655), .B2(new_n688), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1181), .A2(new_n1182), .B1(new_n1185), .B2(new_n916), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1162), .B1(new_n1177), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n932), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1181), .A2(new_n916), .A3(new_n1185), .A4(new_n1182), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT118), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1124), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n717), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1178), .A2(new_n769), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n760), .B1(new_n958), .B2(new_n852), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n787), .A2(new_n343), .B1(new_n1153), .B2(new_n790), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n806), .A2(G125), .B1(new_n795), .B2(G128), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n836), .B2(new_n804), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G132), .C2(new_n798), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT59), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n250), .B(new_n327), .C1(new_n778), .C2(new_n812), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G124), .B2(new_n782), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G97), .A2(new_n798), .B1(new_n806), .B2(G116), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n377), .B2(new_n804), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n779), .A2(G58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n782), .A2(G283), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1053), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n327), .B(new_n287), .C1(new_n794), .C2(new_n531), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1212), .A2(new_n962), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G50), .B1(new_n250), .B2(new_n327), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n467), .B2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1210), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1200), .B1(new_n1222), .B2(new_n772), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1191), .B2(new_n759), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1198), .A2(new_n1226), .ZN(G375));
  OAI21_X1  g1027(.A(new_n760), .B1(G68), .B2(new_n852), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G132), .A2(new_n806), .B1(new_n798), .B2(new_n1154), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n836), .B2(new_n794), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT122), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n467), .B1(new_n787), .B2(new_n348), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n782), .A2(G128), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1213), .B(new_n1235), .C1(new_n812), .C2(new_n790), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(G150), .C2(new_n803), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1232), .A2(new_n1233), .A3(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n799), .A2(new_n247), .B1(new_n531), .B2(new_n804), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1239), .A2(KEYINPUT119), .B1(G294), .B2(new_n806), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(KEYINPUT119), .B2(new_n1239), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT120), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n790), .A2(new_n583), .B1(new_n781), .B2(new_n791), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT121), .Z(new_n1244));
  AOI21_X1  g1044(.A(new_n318), .B1(new_n779), .B2(G77), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n794), .B2(new_n972), .C1(new_n377), .C2(new_n787), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1238), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1228), .B1(new_n1248), .B2(new_n772), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n925), .B2(new_n770), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1130), .B2(new_n758), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT123), .Z(new_n1252));
  NAND2_X1  g1052(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1132), .A2(new_n1010), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT124), .ZN(G381));
  NOR3_X1   g1056(.A1(G396), .A2(G393), .A3(G384), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n753), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1078), .B2(new_n990), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n758), .B1(new_n1259), .B2(new_n1009), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1260), .A2(new_n1261), .B1(new_n984), .B2(new_n980), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1100), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1103), .A2(KEYINPUT115), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1106), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1262), .A3(new_n1266), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1267), .ZN(G407));
  AND3_X1   g1068(.A1(new_n1136), .A2(new_n1140), .A3(new_n1160), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n689), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1198), .A2(new_n1269), .A3(new_n1226), .A4(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT125), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(new_n1273), .A3(G213), .ZN(G409));
  NAND2_X1  g1074(.A1(G390), .A2(new_n1262), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G396), .B(G393), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1266), .ZN(new_n1277));
  AND4_X1   g1077(.A1(KEYINPUT126), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(G387), .B2(new_n1266), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1280), .A2(new_n1276), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1226), .C1(new_n1194), .C2(new_n1197), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT118), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT118), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1010), .B(new_n1193), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1225), .B1(new_n1195), .B2(new_n759), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1269), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1253), .B1(new_n1131), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n717), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1252), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n857), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1252), .A2(G384), .A3(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1290), .A2(new_n1291), .A3(new_n1270), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1271), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1271), .A2(G2897), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1297), .A2(new_n1298), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1301), .B(new_n1302), .C1(new_n1303), .C2(new_n1307), .ZN(new_n1308));
  XOR2_X1   g1108(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1303), .B2(new_n1300), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1282), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1303), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(new_n1299), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1312), .A2(new_n1315), .A3(new_n1317), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1269), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1299), .A3(new_n1283), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1198), .B2(new_n1226), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1283), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1300), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1282), .A2(new_n1322), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1282), .B1(new_n1325), .B2(new_n1322), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


