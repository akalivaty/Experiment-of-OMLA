//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT64), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n223), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n214), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  AOI21_X1  g0047(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT66), .B1(new_n256), .B2(new_n250), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G226), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n251), .A2(KEYINPUT65), .A3(G274), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n249), .B(G274), .C1(G41), .C2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G222), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G223), .A2(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n219), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT67), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n248), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n260), .B(new_n265), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n280), .A2(KEYINPUT70), .A3(G179), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G58), .A2(G68), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n228), .B1(new_n282), .B2(new_n217), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n228), .A2(new_n254), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n254), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n222), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n285), .B1(new_n286), .B2(new_n287), .C1(new_n289), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n227), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n294), .A2(new_n296), .B1(new_n217), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n249), .A2(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G50), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n280), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT70), .B1(new_n280), .B2(G179), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n281), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n299), .B2(new_n302), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n299), .A2(new_n309), .A3(new_n302), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n280), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n280), .A2(KEYINPUT74), .A3(G200), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n315), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n280), .A2(G200), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n313), .A2(new_n317), .A3(new_n318), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n312), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n310), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(new_n315), .A3(KEYINPUT73), .A4(new_n316), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT10), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n308), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n289), .A2(new_n219), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n287), .A2(new_n217), .B1(new_n228), .B2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n296), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n300), .A2(new_n301), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n298), .A2(new_n333), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT12), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n223), .A2(G1698), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n339), .B1(G226), .B2(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n340));
  AND2_X1   g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT75), .B1(new_n340), .B2(new_n342), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n256), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT66), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n248), .A2(new_n251), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G238), .B1(new_n348), .B2(new_n257), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n265), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(new_n350), .A3(KEYINPUT13), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  INV_X1    g0152(.A(new_n265), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n259), .B2(G238), .ZN(new_n354));
  INV_X1    g0154(.A(new_n345), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n248), .A3(new_n343), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G169), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT14), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n346), .B2(new_n350), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n356), .A3(new_n352), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G169), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n360), .A2(new_n361), .A3(G190), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT76), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n338), .B1(new_n363), .B2(G200), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n338), .A2(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n259), .A2(G244), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n269), .A2(G232), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n268), .B(new_n372), .C1(new_n373), .C2(new_n269), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n248), .C1(G107), .C2(new_n268), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n265), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n332), .A2(new_n219), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n297), .A2(G77), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n290), .A2(new_n287), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n228), .A2(new_n219), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT71), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(new_n289), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n378), .B(new_n379), .C1(new_n385), .C2(new_n296), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT72), .ZN(new_n388));
  INV_X1    g0188(.A(new_n376), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G190), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n327), .A2(new_n370), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n275), .B2(new_n228), .ZN(new_n395));
  AND4_X1   g0195(.A1(KEYINPUT7), .A2(new_n266), .A3(new_n228), .A4(new_n267), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n228), .A2(new_n254), .A3(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n282), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n398), .A4(new_n401), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n296), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT78), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n293), .A2(new_n332), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n298), .B2(new_n293), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n404), .A2(new_n405), .A3(new_n410), .A4(new_n296), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n252), .A2(G232), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n265), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n218), .A2(G1698), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n415), .B1(G223), .B2(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n256), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n414), .A2(new_n418), .A3(KEYINPUT79), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  INV_X1    g0220(.A(new_n418), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n252), .A2(G232), .B1(new_n261), .B2(new_n264), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n414), .A2(new_n418), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n424), .A2(new_n304), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT18), .B1(new_n412), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n412), .A2(KEYINPUT18), .A3(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n419), .B2(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n426), .A2(new_n314), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(new_n407), .A3(new_n409), .A4(new_n411), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n389), .A2(new_n425), .ZN(new_n438));
  INV_X1    g0238(.A(new_n386), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n376), .A2(new_n304), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n431), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n394), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n228), .B2(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n213), .A2(KEYINPUT23), .A3(G20), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n254), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n228), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n228), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n268), .A2(new_n456), .A3(new_n228), .A4(G87), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n445), .B1(new_n458), .B2(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n457), .ZN(new_n460));
  INV_X1    g0260(.A(new_n453), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n445), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n296), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n249), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n300), .A2(new_n297), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT25), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n297), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n298), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n470), .A2(G107), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n208), .A2(new_n269), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n268), .B(new_n476), .C1(G257), .C2(new_n269), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n256), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n484), .A2(G264), .A3(new_n256), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(G274), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n481), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n480), .A2(new_n425), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n488), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n479), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(G169), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n475), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(G190), .ZN(new_n495));
  INV_X1    g0295(.A(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n467), .A2(new_n495), .A3(new_n474), .A4(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n298), .A2(new_n450), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n300), .A2(G116), .A3(new_n297), .A4(new_n468), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n295), .A2(new_n227), .B1(G20), .B2(new_n450), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n228), .C1(G33), .C2(new_n209), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n502), .A2(KEYINPUT20), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT20), .B1(new_n502), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n500), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n484), .A2(G270), .A3(new_n256), .ZN(new_n508));
  INV_X1    g0308(.A(G303), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n266), .A2(new_n509), .A3(new_n267), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G264), .A2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n210), .B2(G1698), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n248), .C1(new_n275), .C2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n513), .A3(new_n488), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(G169), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT21), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n507), .A2(new_n514), .A3(new_n517), .A4(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n514), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(G179), .A3(new_n507), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n507), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n514), .A2(new_n314), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(G200), .B2(new_n514), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n373), .A2(new_n269), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n220), .A2(G1698), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n273), .C2(new_n274), .ZN(new_n529));
  INV_X1    g0329(.A(new_n451), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n248), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n487), .A2(new_n248), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n208), .B2(new_n483), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(G200), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n470), .A2(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n384), .A2(new_n298), .ZN(new_n540));
  NOR3_X1   g0340(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n541));
  OR2_X1    g0341(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g0342(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n341), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n228), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n228), .B(G68), .C1(new_n273), .C2(new_n274), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(G97), .A2(new_n288), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n539), .B(new_n540), .C1(new_n549), .C2(new_n300), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n535), .A2(new_n537), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G190), .ZN(new_n554));
  AOI211_X1 g0354(.A(KEYINPUT82), .B(new_n314), .C1(new_n535), .C2(new_n537), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n538), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n287), .A2(new_n219), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  AND2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n564), .B2(G20), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n300), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n469), .A2(new_n209), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n297), .A2(G97), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n208), .B1(new_n266), .B2(new_n267), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(G1698), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(G244), .B1(new_n273), .B2(new_n274), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n572), .B1(G33), .B2(G283), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n572), .A2(G1698), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(G244), .C1(new_n274), .C2(new_n273), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n248), .B1(new_n483), .B2(new_n481), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n578), .A2(new_n248), .B1(G257), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n304), .B1(new_n580), .B2(new_n488), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n220), .B1(new_n266), .B2(new_n267), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n577), .B(new_n503), .C1(new_n582), .C2(KEYINPUT4), .ZN(new_n583));
  OAI21_X1  g0383(.A(G250), .B1(new_n273), .B2(new_n274), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n269), .B1(new_n584), .B2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n248), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(G257), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n488), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n570), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n553), .A2(new_n425), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n540), .B1(new_n384), .B2(new_n469), .C1(new_n549), .C2(new_n300), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n535), .A2(new_n304), .A3(new_n537), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n586), .A2(new_n488), .A3(new_n587), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n586), .A2(G190), .A3(new_n488), .A4(new_n587), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n569), .A3(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n556), .A2(new_n590), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n444), .A2(new_n499), .A3(new_n526), .A4(new_n599), .ZN(G372));
  INV_X1    g0400(.A(new_n430), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n428), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n366), .A2(new_n338), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n441), .B1(new_n369), .B2(new_n368), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n437), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n322), .A2(new_n326), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n308), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n594), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n595), .A2(G169), .ZN(new_n610));
  INV_X1    g0410(.A(new_n567), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n557), .A2(new_n565), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n568), .B1(new_n612), .B2(new_n296), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n610), .A2(new_n588), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n554), .A2(new_n555), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n551), .A2(new_n538), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n594), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n609), .B1(new_n617), .B2(KEYINPUT26), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT86), .B1(new_n581), .B2(new_n589), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n620), .A3(new_n588), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n569), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n535), .A2(G200), .A3(new_n537), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT84), .B1(new_n624), .B2(new_n550), .ZN(new_n625));
  INV_X1    g0425(.A(new_n548), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n544), .A2(new_n228), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n546), .C1(new_n627), .C2(new_n541), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n296), .B1(new_n298), .B2(new_n384), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT84), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n538), .A3(new_n630), .A4(new_n539), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n625), .B(new_n631), .C1(new_n555), .C2(new_n554), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n622), .A2(new_n623), .A3(new_n594), .A4(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n596), .A2(new_n569), .A3(new_n597), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n614), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(new_n498), .A3(new_n594), .A4(new_n632), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n492), .B1(new_n467), .B2(new_n474), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n522), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n519), .A2(KEYINPUT85), .A3(new_n521), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n618), .B(new_n633), .C1(new_n636), .C2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n608), .B1(new_n443), .B2(new_n643), .ZN(G369));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  INV_X1    g0445(.A(G13), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G20), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n249), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  INV_X1    g0450(.A(G213), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(KEYINPUT87), .B(G343), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT88), .Z(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n523), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n645), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n526), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT89), .Z(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n475), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n499), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n494), .B2(new_n655), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n522), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n499), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n637), .A2(new_n655), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT90), .Z(G399));
  NAND2_X1  g0474(.A1(new_n541), .A2(new_n450), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n204), .A2(new_n255), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n231), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n556), .A2(new_n623), .A3(new_n594), .A4(new_n614), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n594), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n631), .B1(new_n555), .B2(new_n554), .ZN(new_n684));
  INV_X1    g0484(.A(new_n625), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n594), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n610), .A2(new_n620), .A3(new_n588), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n620), .B1(new_n610), .B2(new_n588), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n570), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT26), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n494), .A2(KEYINPUT91), .A3(new_n667), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n637), .B2(new_n522), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n683), .B(new_n690), .C1(new_n694), .C2(new_n636), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n655), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(KEYINPUT92), .A3(new_n655), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n642), .A2(new_n655), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n491), .A2(new_n508), .A3(new_n513), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n553), .A3(new_n589), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(KEYINPUT30), .A3(new_n589), .A4(new_n553), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n553), .A2(new_n520), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n425), .A3(new_n496), .A4(new_n595), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n662), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n499), .A2(new_n599), .A3(new_n526), .A4(new_n655), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n703), .B1(G330), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n681), .B1(new_n718), .B2(G1), .ZN(G364));
  NAND2_X1  g0519(.A1(new_n647), .A2(G45), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n677), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n659), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT94), .Z(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n227), .B1(G20), .B2(new_n304), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n425), .A2(new_n432), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n228), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n333), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n228), .B1(new_n733), .B2(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n209), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n425), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n275), .B(new_n735), .C1(G77), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n432), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G107), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n730), .A2(new_n733), .ZN(new_n744));
  INV_X1    g0544(.A(G159), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT32), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n228), .A2(new_n314), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n740), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n207), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n729), .A2(new_n748), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(G50), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n739), .A2(new_n743), .A3(new_n747), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n748), .A2(new_n736), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n732), .B(new_n754), .C1(G58), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n731), .ZN(new_n758));
  INV_X1    g0558(.A(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n744), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G329), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n742), .A2(G283), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G326), .B2(new_n752), .ZN(new_n767));
  INV_X1    g0567(.A(new_n749), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G303), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n268), .B1(new_n756), .B2(G322), .ZN(new_n770));
  INV_X1    g0570(.A(new_n734), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G294), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n767), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G311), .B2(new_n738), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n728), .B1(new_n757), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n275), .A2(new_n204), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n231), .A2(new_n482), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n482), .C2(new_n243), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n268), .A2(new_n204), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(G116), .B2(new_n204), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n725), .A2(new_n728), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n727), .A2(new_n775), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G330), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n722), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n660), .A3(new_n721), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(G396));
  NOR2_X1   g0589(.A1(new_n441), .A2(new_n662), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n662), .A2(new_n439), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n393), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(new_n441), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n701), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n642), .A2(new_n655), .A3(new_n793), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n717), .A2(G330), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n797), .B(new_n798), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n721), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n793), .A2(new_n724), .ZN(new_n801));
  INV_X1    g0601(.A(new_n728), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n756), .B1(new_n738), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n751), .C1(new_n286), .C2(new_n731), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT34), .Z(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G50), .B2(new_n768), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n275), .B1(new_n763), .B2(G132), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n771), .A2(G58), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n741), .A2(new_n333), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n735), .B1(G311), .B2(new_n763), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n213), .B2(new_n749), .ZN(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n275), .B1(new_n755), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n742), .A2(G87), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n450), .B2(new_n737), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT95), .B(G283), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(new_n509), .B2(new_n751), .C1(new_n731), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n802), .B1(new_n812), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n801), .A2(new_n721), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n728), .A2(new_n723), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(G77), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n800), .A2(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n412), .A2(new_n427), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n412), .A2(new_n652), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n831), .A3(new_n436), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n431), .B2(new_n437), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n406), .A2(new_n409), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n652), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT97), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(new_n840), .A3(new_n652), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT17), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n436), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n602), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n427), .A2(new_n837), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n436), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n436), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n836), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n716), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n711), .A2(KEYINPUT99), .A3(KEYINPUT31), .A4(new_n662), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(new_n714), .A3(new_n715), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n793), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n662), .A2(new_n338), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n366), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n370), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n861), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n848), .A2(new_n849), .ZN(new_n865));
  INV_X1    g0665(.A(new_n842), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n431), .B2(new_n437), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n829), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n851), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n863), .A2(KEYINPUT40), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n444), .A2(new_n856), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(G330), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT98), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n703), .B2(new_n444), .ZN(new_n875));
  AOI211_X1 g0675(.A(KEYINPUT98), .B(new_n443), .C1(new_n700), .C2(new_n702), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(new_n608), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n873), .B(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n603), .A2(new_n662), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n431), .A2(new_n652), .ZN(new_n885));
  INV_X1    g0685(.A(new_n790), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n861), .B1(new_n796), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n879), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n249), .B2(new_n647), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n564), .B(KEYINPUT96), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n450), .B1(new_n892), .B2(KEYINPUT35), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(new_n229), .C1(KEYINPUT35), .C2(new_n892), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n231), .A2(G77), .A3(new_n399), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(G50), .B2(new_n333), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G1), .A3(new_n646), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n891), .A2(new_n895), .A3(new_n898), .ZN(G367));
  NAND2_X1  g0699(.A1(new_n662), .A2(new_n550), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT100), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n609), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT101), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n901), .B2(new_n686), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT43), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n635), .B1(new_n569), .B2(new_n655), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n622), .A2(new_n662), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n637), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n662), .B1(new_n913), .B2(new_n590), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n499), .A2(new_n635), .A3(new_n668), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n908), .B1(new_n909), .B2(new_n906), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n908), .A2(new_n914), .A3(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n666), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n912), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n677), .B(KEYINPUT41), .Z(new_n923));
  INV_X1    g0723(.A(KEYINPUT104), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n672), .B2(new_n912), .ZN(new_n926));
  INV_X1    g0726(.A(new_n912), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n671), .A2(new_n927), .A3(KEYINPUT103), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT45), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n671), .A2(new_n927), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT44), .Z(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n926), .B2(new_n928), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n920), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n666), .A2(new_n932), .A3(new_n933), .A4(new_n930), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n924), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n669), .B1(new_n665), .B2(new_n668), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n660), .B(new_n939), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n718), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n937), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n718), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n923), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n720), .A2(G1), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n922), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n906), .A2(new_n726), .ZN(new_n948));
  INV_X1    g0748(.A(new_n721), .ZN(new_n949));
  INV_X1    g0749(.A(new_n777), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n783), .B1(new_n204), .B2(new_n384), .C1(new_n239), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n742), .A2(G97), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n749), .A2(new_n450), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(KEYINPUT46), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n268), .B1(new_n953), .B2(KEYINPUT46), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n213), .B2(new_n734), .C1(new_n815), .C2(new_n731), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(new_n738), .C2(new_n820), .ZN(new_n957));
  XNOR2_X1  g0757(.A(KEYINPUT105), .B(G311), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n751), .A2(new_n958), .B1(new_n755), .B2(new_n509), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT106), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(new_n759), .C2(new_n744), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n742), .A2(G77), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n217), .B2(new_n737), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G150), .A2(new_n756), .B1(new_n763), .B2(G137), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n333), .B2(new_n734), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G58), .C2(new_n768), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n752), .A2(G143), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n758), .A2(G159), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n966), .A2(new_n268), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  OAI211_X1 g0771(.A(new_n949), .B(new_n951), .C1(new_n971), .C2(new_n802), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n948), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n947), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(G387));
  OAI211_X1 g0775(.A(new_n664), .B(new_n726), .C1(new_n494), .C2(new_n655), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n236), .A2(G45), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n290), .A2(G50), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT108), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT50), .Z(new_n981));
  AOI21_X1  g0781(.A(G45), .B1(G68), .B2(G77), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n676), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n777), .A3(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(G107), .B2(new_n204), .C1(new_n676), .C2(new_n781), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n783), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n384), .A2(new_n734), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G150), .B2(new_n763), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n952), .C1(new_n217), .C2(new_n755), .ZN(new_n989));
  INV_X1    g0789(.A(new_n293), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n990), .A2(new_n758), .B1(G77), .B2(new_n768), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n333), .B2(new_n737), .C1(new_n745), .C2(new_n751), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n989), .A2(new_n992), .A3(new_n275), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G322), .A2(new_n752), .B1(new_n756), .B2(G317), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n509), .B2(new_n737), .C1(new_n731), .C2(new_n958), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT48), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n815), .B2(new_n749), .C1(new_n734), .C2(new_n821), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT49), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n741), .A2(new_n450), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n268), .B(new_n999), .C1(G326), .C2(new_n763), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n993), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n986), .B(new_n949), .C1(new_n1001), .C2(new_n802), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT109), .Z(new_n1003));
  AOI22_X1  g0803(.A1(new_n940), .A2(new_n945), .B1(new_n976), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n677), .B(KEYINPUT110), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n941), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n940), .A2(new_n718), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G393));
  INV_X1    g0809(.A(new_n942), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n935), .A2(new_n936), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1005), .B1(new_n1011), .B2(new_n941), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n935), .A2(new_n936), .A3(new_n945), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G317), .A2(new_n752), .B1(new_n756), .B2(G311), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT52), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G116), .B2(new_n771), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n743), .B1(new_n815), .B2(new_n737), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n268), .B(new_n1018), .C1(G322), .C2(new_n763), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n509), .B2(new_n731), .C1(new_n749), .C2(new_n821), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n734), .A2(new_n219), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n768), .A2(G68), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n737), .B2(new_n290), .C1(new_n217), .C2(new_n731), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G143), .C2(new_n763), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n751), .A2(new_n286), .B1(new_n755), .B2(new_n745), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n268), .A3(new_n817), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n802), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n783), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n204), .A2(new_n209), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n777), .C2(new_n246), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1029), .A2(new_n721), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n725), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n912), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1013), .A2(new_n1014), .A3(new_n1035), .ZN(G390));
  AOI21_X1  g0836(.A(new_n882), .B1(new_n836), .B2(new_n851), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n698), .A2(new_n699), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n792), .A2(new_n441), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n790), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1040), .B2(new_n861), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n796), .A2(new_n886), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n370), .A2(new_n858), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n860), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n882), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(KEYINPUT111), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n887), .B2(new_n882), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT39), .B1(new_n836), .B2(new_n851), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1048), .B(new_n1050), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1045), .A2(new_n717), .A3(G330), .A4(new_n793), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1041), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT111), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n887), .A2(new_n1049), .A3(new_n882), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n881), .A2(new_n883), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n698), .A2(new_n699), .B1(new_n441), .B2(new_n792), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1045), .B1(new_n1060), .B2(new_n790), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1058), .A2(new_n1059), .B1(new_n1061), .B2(new_n1037), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n862), .A2(G330), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n945), .B(new_n1055), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1059), .A2(new_n723), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n741), .A2(new_n217), .B1(new_n734), .B2(new_n745), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n731), .A2(new_n804), .B1(new_n737), .B2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1066), .B(new_n1069), .C1(G132), .C2(new_n756), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n763), .A2(G125), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n749), .A2(new_n286), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT53), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n275), .B1(new_n752), .B2(G128), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n275), .B1(new_n731), .B2(new_n213), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1076), .A2(new_n750), .A3(new_n810), .A4(new_n1022), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n756), .A2(G116), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n752), .A2(G283), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G97), .A2(new_n738), .B1(new_n763), .B2(G294), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n802), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n721), .B(new_n1082), .C1(new_n293), .C2(new_n825), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT114), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n1065), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1064), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1064), .A2(KEYINPUT115), .A3(new_n1085), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n871), .A2(G330), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n608), .C1(new_n875), .C2(new_n876), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n861), .B1(new_n798), .B2(new_n794), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1063), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1042), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n861), .B1(new_n857), .B2(new_n786), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1040), .A2(new_n1054), .A3(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT112), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1063), .B1(new_n1041), .B2(new_n1053), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n877), .A2(new_n608), .A3(new_n1092), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT112), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1103), .A2(new_n1107), .A3(new_n1006), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1090), .A2(new_n1091), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1091), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G378));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1093), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1106), .B2(new_n1099), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n863), .A2(KEYINPUT40), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n864), .A2(new_n869), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n786), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n889), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n884), .B(new_n888), .C1(new_n870), .C2(new_n786), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n327), .B(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n303), .A2(new_n652), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1122), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1120), .A2(new_n1121), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1113), .B1(new_n1116), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1120), .A2(new_n1121), .A3(new_n1130), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(KEYINPUT57), .A3(new_n1115), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1135), .A2(new_n1006), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n723), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G41), .B1(new_n763), .B2(G124), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n756), .A2(G128), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G132), .A2(new_n758), .B1(new_n738), .B2(G137), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G125), .C2(new_n752), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n286), .B2(new_n734), .C1(new_n749), .C2(new_n1067), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n254), .B(new_n1142), .C1(new_n1147), .C2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n745), .B2(new_n741), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT58), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n255), .B1(new_n734), .B2(new_n333), .C1(new_n219), .C2(new_n749), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n758), .A2(G97), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n742), .A2(G58), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n763), .A2(G283), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n275), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G116), .C2(new_n752), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n213), .B2(new_n755), .C1(new_n384), .C2(new_n737), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1150), .A2(new_n1151), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1152), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n217), .B1(new_n273), .B2(G41), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT117), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT118), .Z(new_n1166));
  OAI21_X1  g0966(.A(new_n728), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n825), .A2(new_n217), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1141), .A2(new_n949), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT121), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n945), .B2(new_n1138), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1140), .A2(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1105), .A2(new_n923), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n826), .A2(G68), .ZN(new_n1176));
  INV_X1    g0976(.A(G132), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n268), .B1(new_n751), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G159), .A2(new_n768), .B1(new_n742), .B2(G58), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n804), .B2(new_n755), .C1(new_n731), .C2(new_n1067), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G128), .C2(new_n763), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n217), .B2(new_n734), .C1(new_n286), .C2(new_n737), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n737), .A2(new_n213), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1183), .B(new_n987), .C1(G116), .C2(new_n758), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n268), .B1(new_n756), .B2(G283), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n749), .A2(new_n209), .B1(new_n744), .B2(new_n509), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT123), .Z(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n962), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n751), .A2(new_n815), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT124), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n721), .B(new_n1176), .C1(new_n1191), .C2(new_n728), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n861), .A2(new_n723), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT122), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1104), .A2(new_n945), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1175), .A2(new_n1195), .ZN(G381));
  INV_X1    g0996(.A(G390), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n974), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1198), .A2(G396), .A3(G393), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G381), .A2(G384), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1090), .A2(new_n1108), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G375), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(G407));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  OAI211_X1 g1004(.A(G407), .B(G213), .C1(new_n653), .C2(new_n1204), .ZN(G409));
  INV_X1    g1005(.A(KEYINPUT126), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n653), .A2(new_n651), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT60), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1174), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1093), .A2(new_n1099), .A3(KEYINPUT60), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1006), .A3(new_n1105), .A4(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(G384), .A3(new_n1195), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G384), .B1(new_n1211), .B2(new_n1195), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G2897), .B(new_n1207), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1207), .A2(G2897), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1212), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1201), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1169), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1115), .A2(new_n923), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1134), .B1(new_n1222), .B2(new_n946), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1220), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1111), .B2(G375), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1207), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1206), .B1(new_n1227), .B2(KEYINPUT61), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1172), .B(new_n1140), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1207), .B1(new_n1230), .B2(new_n1224), .ZN(new_n1231));
  OAI211_X1 g1031(.A(KEYINPUT126), .B(new_n1229), .C1(new_n1231), .C2(new_n1219), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1236), .A3(new_n1233), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1228), .A2(new_n1232), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT125), .B1(new_n974), .B2(new_n1197), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(G396), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G390), .B1(new_n947), .B2(new_n973), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1238), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1234), .B1(new_n1227), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1233), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n1229), .A3(new_n1244), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(G405));
  NAND2_X1  g1051(.A1(new_n1233), .A2(KEYINPUT127), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1240), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1233), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(new_n1220), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1230), .B2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1260), .B(new_n1263), .ZN(G402));
endmodule


