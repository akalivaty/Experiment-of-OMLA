

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761;

  OR2_X1 U371 ( .A1(n527), .A2(n526), .ZN(n540) );
  NOR2_X1 U372 ( .A1(n529), .A2(n528), .ZN(n652) );
  INV_X1 U373 ( .A(G953), .ZN(n754) );
  NOR2_X1 U374 ( .A1(n699), .A2(n529), .ZN(n524) );
  XNOR2_X2 U375 ( .A(n623), .B(n622), .ZN(n735) );
  XNOR2_X2 U376 ( .A(n408), .B(n407), .ZN(n500) );
  XNOR2_X1 U377 ( .A(n604), .B(n603), .ZN(n621) );
  XNOR2_X1 U378 ( .A(n413), .B(n351), .ZN(n594) );
  NAND2_X1 U379 ( .A1(n621), .A2(n424), .ZN(n623) );
  AND2_X1 U380 ( .A1(n633), .A2(n632), .ZN(n602) );
  XNOR2_X1 U381 ( .A(n587), .B(n586), .ZN(n633) );
  AND2_X1 U382 ( .A1(n568), .A2(n669), .ZN(n570) );
  BUF_X1 U383 ( .A(n594), .Z(n595) );
  OR2_X1 U384 ( .A1(n730), .A2(G902), .ZN(n413) );
  OR2_X1 U385 ( .A1(n716), .A2(n485), .ZN(n490) );
  XNOR2_X1 U386 ( .A(n479), .B(n478), .ZN(n740) );
  XNOR2_X1 U387 ( .A(n741), .B(KEYINPUT70), .ZN(n477) );
  XNOR2_X1 U388 ( .A(n392), .B(n391), .ZN(n741) );
  XNOR2_X1 U389 ( .A(n462), .B(n461), .ZN(n479) );
  XNOR2_X1 U390 ( .A(n446), .B(G128), .ZN(n408) );
  XNOR2_X1 U391 ( .A(n450), .B(G110), .ZN(n392) );
  XOR2_X1 U392 ( .A(KEYINPUT3), .B(G119), .Z(n461) );
  INV_X1 U393 ( .A(KEYINPUT65), .ZN(n446) );
  XNOR2_X1 U394 ( .A(KEYINPUT77), .B(G143), .ZN(n407) );
  XNOR2_X1 U395 ( .A(G116), .B(G113), .ZN(n460) );
  XNOR2_X1 U396 ( .A(KEYINPUT16), .B(G122), .ZN(n478) );
  XNOR2_X1 U397 ( .A(G101), .B(KEYINPUT72), .ZN(n450) );
  XNOR2_X1 U398 ( .A(G107), .B(G104), .ZN(n391) );
  NOR2_X2 U399 ( .A1(n735), .A2(n752), .ZN(n349) );
  INV_X1 U400 ( .A(n692), .ZN(n350) );
  NOR2_X1 U401 ( .A1(n735), .A2(n752), .ZN(n625) );
  XNOR2_X1 U402 ( .A(n571), .B(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U403 ( .A1(n559), .A2(n517), .ZN(n518) );
  XNOR2_X1 U404 ( .A(n484), .B(n370), .ZN(n369) );
  XNOR2_X1 U405 ( .A(n740), .B(n477), .ZN(n372) );
  XNOR2_X1 U406 ( .A(n481), .B(n371), .ZN(n370) );
  INV_X1 U407 ( .A(n729), .ZN(n381) );
  INV_X1 U408 ( .A(G237), .ZN(n458) );
  OR2_X1 U409 ( .A1(n659), .A2(n644), .ZN(n614) );
  XOR2_X1 U410 ( .A(G125), .B(G146), .Z(n482) );
  XNOR2_X1 U411 ( .A(n527), .B(KEYINPUT38), .ZN(n683) );
  XNOR2_X1 U412 ( .A(n501), .B(n365), .ZN(n553) );
  XNOR2_X1 U413 ( .A(n366), .B(G478), .ZN(n365) );
  INV_X1 U414 ( .A(KEYINPUT100), .ZN(n366) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n448) );
  NAND2_X1 U416 ( .A1(n395), .A2(n393), .ZN(n752) );
  AND2_X1 U417 ( .A1(n758), .A2(n394), .ZN(n393) );
  XNOR2_X1 U418 ( .A(n397), .B(n396), .ZN(n395) );
  INV_X1 U419 ( .A(n665), .ZN(n394) );
  XNOR2_X1 U420 ( .A(G140), .B(G137), .ZN(n449) );
  XNOR2_X1 U421 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n425) );
  XNOR2_X1 U422 ( .A(n482), .B(n368), .ZN(n746) );
  INV_X1 U423 ( .A(KEYINPUT10), .ZN(n368) );
  XNOR2_X1 U424 ( .A(G119), .B(G128), .ZN(n427) );
  XNOR2_X1 U425 ( .A(n495), .B(n494), .ZN(n367) );
  XNOR2_X1 U426 ( .A(G116), .B(G107), .ZN(n493) );
  XNOR2_X1 U427 ( .A(n607), .B(n606), .ZN(n678) );
  INV_X1 U428 ( .A(KEYINPUT0), .ZN(n414) );
  BUF_X1 U429 ( .A(n568), .Z(n670) );
  AND2_X1 U430 ( .A1(n384), .A2(n389), .ZN(n383) );
  NAND2_X1 U431 ( .A1(n729), .A2(n387), .ZN(n386) );
  NAND2_X1 U432 ( .A1(n718), .A2(n385), .ZN(n384) );
  AND2_X1 U433 ( .A1(n378), .A2(KEYINPUT56), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n354), .B(n482), .ZN(n371) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U437 ( .A(G143), .B(G140), .ZN(n507) );
  XOR2_X1 U438 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n508) );
  XNOR2_X1 U439 ( .A(G113), .B(G131), .ZN(n505) );
  NAND2_X1 U440 ( .A1(n364), .A2(n704), .ZN(n416) );
  NAND2_X1 U441 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n440) );
  XOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT71), .Z(n464) );
  XNOR2_X1 U444 ( .A(G101), .B(G146), .ZN(n465) );
  XOR2_X1 U445 ( .A(KEYINPUT92), .B(G137), .Z(n466) );
  INV_X1 U446 ( .A(G210), .ZN(n385) );
  AND2_X1 U447 ( .A1(n390), .A2(G210), .ZN(n387) );
  NAND2_X1 U448 ( .A1(n405), .A2(n406), .ZN(n404) );
  NAND2_X1 U449 ( .A1(n588), .A2(n682), .ZN(n405) );
  XNOR2_X1 U450 ( .A(n492), .B(n491), .ZN(n559) );
  XNOR2_X1 U451 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U452 ( .A(n746), .B(n425), .ZN(n431) );
  XNOR2_X1 U453 ( .A(n353), .B(n367), .ZN(n498) );
  XNOR2_X1 U454 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U455 ( .A(n747), .B(n352), .ZN(n374) );
  XNOR2_X1 U456 ( .A(KEYINPUT74), .B(G146), .ZN(n452) );
  XNOR2_X1 U457 ( .A(n567), .B(n566), .ZN(n758) );
  XNOR2_X1 U458 ( .A(n601), .B(n600), .ZN(n642) );
  AND2_X1 U459 ( .A1(n423), .A2(n598), .ZN(n421) );
  XNOR2_X1 U460 ( .A(n610), .B(n609), .ZN(n659) );
  XNOR2_X1 U461 ( .A(KEYINPUT101), .B(n516), .ZN(n656) );
  NAND2_X1 U462 ( .A1(n379), .A2(n377), .ZN(n376) );
  XNOR2_X1 U463 ( .A(n436), .B(n435), .ZN(n351) );
  XOR2_X1 U464 ( .A(n477), .B(n453), .Z(n352) );
  XOR2_X1 U465 ( .A(n493), .B(KEYINPUT99), .Z(n353) );
  XOR2_X1 U466 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n354) );
  XNOR2_X1 U467 ( .A(n593), .B(n592), .ZN(n599) );
  AND2_X1 U468 ( .A1(n599), .A2(n598), .ZN(n355) );
  XOR2_X1 U469 ( .A(n590), .B(KEYINPUT103), .Z(n356) );
  AND2_X1 U470 ( .A1(n402), .A2(n400), .ZN(n357) );
  AND2_X1 U471 ( .A1(n375), .A2(n380), .ZN(n358) );
  NAND2_X1 U472 ( .A1(n349), .A2(KEYINPUT2), .ZN(n359) );
  AND2_X1 U473 ( .A1(n612), .A2(n542), .ZN(n360) );
  INV_X1 U474 ( .A(KEYINPUT41), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n372), .B(n369), .ZN(n716) );
  AND2_X1 U476 ( .A1(n682), .A2(KEYINPUT41), .ZN(n361) );
  AND2_X1 U477 ( .A1(n718), .A2(n388), .ZN(n362) );
  XOR2_X1 U478 ( .A(n627), .B(n626), .Z(n363) );
  INV_X1 U479 ( .A(n734), .ZN(n389) );
  INV_X1 U480 ( .A(KEYINPUT56), .ZN(n388) );
  NAND2_X1 U481 ( .A1(n374), .A2(n459), .ZN(n412) );
  NAND2_X1 U482 ( .A1(n625), .A2(KEYINPUT82), .ZN(n364) );
  NAND2_X1 U483 ( .A1(n415), .A2(n418), .ZN(n417) );
  AND2_X1 U484 ( .A1(n588), .A2(n361), .ZN(n403) );
  XNOR2_X1 U485 ( .A(n432), .B(n433), .ZN(n730) );
  AND2_X1 U486 ( .A1(n409), .A2(n542), .ZN(n457) );
  NAND2_X1 U487 ( .A1(n401), .A2(n406), .ZN(n400) );
  XNOR2_X1 U488 ( .A(n542), .B(KEYINPUT1), .ZN(n568) );
  NAND2_X1 U489 ( .A1(n570), .A2(n373), .ZN(n607) );
  INV_X1 U490 ( .A(n605), .ZN(n373) );
  XNOR2_X1 U491 ( .A(n374), .B(n721), .ZN(n722) );
  NAND2_X1 U492 ( .A1(n382), .A2(n388), .ZN(n375) );
  NAND2_X1 U493 ( .A1(n386), .A2(n383), .ZN(n382) );
  NAND2_X1 U494 ( .A1(n358), .A2(n376), .ZN(G51) );
  NAND2_X1 U495 ( .A1(n381), .A2(n718), .ZN(n378) );
  INV_X1 U496 ( .A(n382), .ZN(n379) );
  NAND2_X1 U497 ( .A1(n381), .A2(n362), .ZN(n380) );
  INV_X1 U498 ( .A(n718), .ZN(n390) );
  NOR2_X2 U499 ( .A1(n476), .A2(n475), .ZN(n555) );
  NAND2_X1 U500 ( .A1(n398), .A2(n550), .ZN(n397) );
  AND2_X1 U501 ( .A1(n551), .A2(n399), .ZN(n398) );
  INV_X1 U502 ( .A(n651), .ZN(n399) );
  NAND2_X1 U503 ( .A1(n404), .A2(n357), .ZN(n699) );
  INV_X1 U504 ( .A(n683), .ZN(n401) );
  NAND2_X1 U505 ( .A1(n403), .A2(n683), .ZN(n402) );
  NAND2_X1 U506 ( .A1(n683), .A2(n682), .ZN(n687) );
  XNOR2_X2 U507 ( .A(n483), .B(n448), .ZN(n471) );
  XNOR2_X2 U508 ( .A(n500), .B(n447), .ZN(n483) );
  OR2_X1 U509 ( .A1(n594), .A2(n666), .ZN(n611) );
  NOR2_X1 U510 ( .A1(n594), .A2(n410), .ZN(n409) );
  NAND2_X1 U511 ( .A1(n411), .A2(n589), .ZN(n410) );
  INV_X1 U512 ( .A(n520), .ZN(n411) );
  XNOR2_X2 U513 ( .A(n412), .B(n456), .ZN(n542) );
  NAND2_X1 U514 ( .A1(n608), .A2(n356), .ZN(n593) );
  NAND2_X1 U515 ( .A1(n608), .A2(n360), .ZN(n613) );
  XNOR2_X2 U516 ( .A(n580), .B(n414), .ZN(n608) );
  NAND2_X1 U517 ( .A1(n416), .A2(n485), .ZN(n415) );
  AND2_X4 U518 ( .A1(n417), .A2(n359), .ZN(n729) );
  INV_X1 U519 ( .A(KEYINPUT82), .ZN(n419) );
  NAND2_X1 U520 ( .A1(n349), .A2(n485), .ZN(n420) );
  NAND2_X1 U521 ( .A1(n599), .A2(n421), .ZN(n601) );
  NAND2_X1 U522 ( .A1(n355), .A2(n618), .ZN(n619) );
  BUF_X1 U523 ( .A(n729), .Z(n725) );
  XOR2_X1 U524 ( .A(n428), .B(n427), .Z(n422) );
  AND2_X1 U525 ( .A1(n670), .A2(n595), .ZN(n423) );
  AND2_X1 U526 ( .A1(n620), .A2(n759), .ZN(n424) );
  INV_X1 U527 ( .A(n611), .ZN(n669) );
  INV_X1 U528 ( .A(KEYINPUT44), .ZN(n603) );
  XNOR2_X1 U529 ( .A(n460), .B(KEYINPUT69), .ZN(n462) );
  XNOR2_X1 U530 ( .A(n730), .B(KEYINPUT124), .ZN(n731) );
  XNOR2_X1 U531 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U532 ( .A(n449), .B(KEYINPUT90), .Z(n433) );
  NAND2_X1 U533 ( .A1(G234), .A2(n754), .ZN(n426) );
  XOR2_X1 U534 ( .A(KEYINPUT8), .B(n426), .Z(n496) );
  NAND2_X1 U535 ( .A1(G221), .A2(n496), .ZN(n429) );
  XOR2_X1 U536 ( .A(KEYINPUT81), .B(G110), .Z(n428) );
  XNOR2_X1 U537 ( .A(n429), .B(n422), .ZN(n430) );
  XNOR2_X1 U538 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U539 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n436) );
  XNOR2_X1 U540 ( .A(KEYINPUT15), .B(G902), .ZN(n624) );
  NAND2_X1 U541 ( .A1(n624), .A2(G234), .ZN(n434) );
  XNOR2_X1 U542 ( .A(n434), .B(KEYINPUT20), .ZN(n437) );
  NAND2_X1 U543 ( .A1(n437), .A2(G217), .ZN(n435) );
  NAND2_X1 U544 ( .A1(n437), .A2(G221), .ZN(n439) );
  INV_X1 U545 ( .A(KEYINPUT21), .ZN(n438) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n589) );
  INV_X1 U547 ( .A(n589), .ZN(n666) );
  XNOR2_X1 U548 ( .A(n440), .B(KEYINPUT14), .ZN(n442) );
  NAND2_X1 U549 ( .A1(G952), .A2(n442), .ZN(n441) );
  XNOR2_X1 U550 ( .A(KEYINPUT88), .B(n441), .ZN(n698) );
  NOR2_X1 U551 ( .A1(G953), .A2(n698), .ZN(n575) );
  NAND2_X1 U552 ( .A1(G902), .A2(n442), .ZN(n572) );
  NOR2_X1 U553 ( .A1(G900), .A2(n572), .ZN(n443) );
  NAND2_X1 U554 ( .A1(G953), .A2(n443), .ZN(n444) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(n444), .Z(n445) );
  NOR2_X1 U556 ( .A1(n575), .A2(n445), .ZN(n520) );
  XNOR2_X1 U557 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n447) );
  XNOR2_X2 U558 ( .A(n471), .B(n449), .ZN(n747) );
  NAND2_X1 U559 ( .A1(n754), .A2(G227), .ZN(n451) );
  XNOR2_X1 U560 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U561 ( .A(KEYINPUT68), .B(G469), .ZN(n455) );
  INV_X1 U562 ( .A(KEYINPUT67), .ZN(n454) );
  XNOR2_X1 U563 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n457), .B(KEYINPUT73), .ZN(n476) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n474) );
  INV_X1 U566 ( .A(G902), .ZN(n459) );
  NAND2_X1 U567 ( .A1(n459), .A2(n458), .ZN(n486) );
  NAND2_X1 U568 ( .A1(n486), .A2(G214), .ZN(n682) );
  NAND2_X1 U569 ( .A1(n502), .A2(G210), .ZN(n463) );
  XNOR2_X1 U570 ( .A(n464), .B(n463), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n479), .B(n469), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n627) );
  OR2_X1 U575 ( .A1(n627), .A2(G902), .ZN(n472) );
  XNOR2_X2 U576 ( .A(n472), .B(G472), .ZN(n676) );
  NAND2_X1 U577 ( .A1(n682), .A2(n676), .ZN(n473) );
  XOR2_X1 U578 ( .A(n474), .B(n473), .Z(n475) );
  NAND2_X1 U579 ( .A1(n754), .A2(G224), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n480), .B(KEYINPUT86), .ZN(n481) );
  INV_X1 U581 ( .A(n483), .ZN(n484) );
  INV_X1 U582 ( .A(n624), .ZN(n485) );
  NAND2_X1 U583 ( .A1(n486), .A2(G210), .ZN(n488) );
  INV_X1 U584 ( .A(KEYINPUT87), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X2 U586 ( .A(n490), .B(n489), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n555), .A2(n683), .ZN(n492) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n495) );
  XNOR2_X1 U589 ( .A(G134), .B(G122), .ZN(n494) );
  NAND2_X1 U590 ( .A1(G217), .A2(n496), .ZN(n497) );
  XNOR2_X1 U591 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n500), .B(n499), .ZN(n726) );
  NOR2_X1 U593 ( .A1(n726), .A2(G902), .ZN(n501) );
  INV_X1 U594 ( .A(n553), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  XOR2_X1 U596 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n504) );
  NAND2_X1 U597 ( .A1(G214), .A2(n502), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n504), .B(n503), .ZN(n512) );
  XOR2_X1 U599 ( .A(G122), .B(G104), .Z(n506) );
  XNOR2_X1 U600 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U601 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U602 ( .A(n510), .B(n509), .Z(n511) );
  XNOR2_X1 U603 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n746), .B(n513), .ZN(n636) );
  NOR2_X1 U605 ( .A1(G902), .A2(n636), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n530), .A2(n552), .ZN(n516) );
  INV_X1 U608 ( .A(n656), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n518), .B(KEYINPUT40), .ZN(n761) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n588) );
  INV_X1 U611 ( .A(n588), .ZN(n685) );
  XOR2_X1 U612 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n522) );
  NAND2_X1 U613 ( .A1(n594), .A2(n589), .ZN(n519) );
  NOR2_X1 U614 ( .A1(n520), .A2(n519), .ZN(n537) );
  NAND2_X1 U615 ( .A1(n373), .A2(n537), .ZN(n521) );
  XNOR2_X1 U616 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U617 ( .A1(n523), .A2(n542), .ZN(n529) );
  XNOR2_X1 U618 ( .A(n524), .B(KEYINPUT42), .ZN(n760) );
  NOR2_X1 U619 ( .A1(n761), .A2(n760), .ZN(n525) );
  XNOR2_X1 U620 ( .A(n525), .B(KEYINPUT46), .ZN(n551) );
  INV_X1 U621 ( .A(n682), .ZN(n526) );
  XNOR2_X2 U622 ( .A(n540), .B(KEYINPUT19), .ZN(n579) );
  INV_X1 U623 ( .A(n579), .ZN(n528) );
  NOR2_X1 U624 ( .A1(n552), .A2(n530), .ZN(n531) );
  XNOR2_X1 U625 ( .A(KEYINPUT102), .B(n531), .ZN(n660) );
  NOR2_X1 U626 ( .A1(n660), .A2(n656), .ZN(n688) );
  INV_X1 U627 ( .A(n688), .ZN(n615) );
  NAND2_X1 U628 ( .A1(n652), .A2(n615), .ZN(n532) );
  INV_X1 U629 ( .A(KEYINPUT47), .ZN(n533) );
  NAND2_X1 U630 ( .A1(n532), .A2(n533), .ZN(n536) );
  NAND2_X1 U631 ( .A1(KEYINPUT80), .A2(n533), .ZN(n534) );
  NAND2_X1 U632 ( .A1(n652), .A2(n534), .ZN(n535) );
  NAND2_X1 U633 ( .A1(n536), .A2(n535), .ZN(n544) );
  INV_X1 U634 ( .A(n537), .ZN(n538) );
  XNOR2_X1 U635 ( .A(n676), .B(KEYINPUT6), .ZN(n598) );
  NOR2_X1 U636 ( .A1(n538), .A2(n598), .ZN(n539) );
  NAND2_X1 U637 ( .A1(n656), .A2(n539), .ZN(n561) );
  NOR2_X1 U638 ( .A1(n561), .A2(n540), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n541), .B(KEYINPUT36), .ZN(n543) );
  NAND2_X1 U640 ( .A1(n543), .A2(n670), .ZN(n663) );
  NAND2_X1 U641 ( .A1(n544), .A2(n663), .ZN(n549) );
  INV_X1 U642 ( .A(n652), .ZN(n545) );
  NOR2_X1 U643 ( .A1(n545), .A2(KEYINPUT80), .ZN(n546) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(n546), .ZN(n547) );
  NOR2_X1 U645 ( .A1(n547), .A2(n615), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n549), .A2(n548), .ZN(n550) );
  AND2_X1 U647 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U648 ( .A(n554), .B(KEYINPUT105), .ZN(n583) );
  INV_X1 U649 ( .A(n527), .ZN(n556) );
  NAND2_X1 U650 ( .A1(n555), .A2(n556), .ZN(n557) );
  XOR2_X1 U651 ( .A(KEYINPUT109), .B(n557), .Z(n558) );
  NOR2_X1 U652 ( .A1(n583), .A2(n558), .ZN(n651) );
  INV_X1 U653 ( .A(n660), .ZN(n560) );
  NOR2_X1 U654 ( .A1(n560), .A2(n559), .ZN(n665) );
  INV_X1 U655 ( .A(n561), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n682), .A2(n562), .ZN(n563) );
  OR2_X1 U657 ( .A1(n670), .A2(n563), .ZN(n564) );
  XNOR2_X1 U658 ( .A(n564), .B(KEYINPUT43), .ZN(n565) );
  NAND2_X1 U659 ( .A1(n565), .A2(n527), .ZN(n567) );
  INV_X1 U660 ( .A(KEYINPUT107), .ZN(n566) );
  INV_X1 U661 ( .A(n598), .ZN(n569) );
  NAND2_X1 U662 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U663 ( .A(n572), .ZN(n573) );
  NOR2_X1 U664 ( .A1(G898), .A2(n754), .ZN(n742) );
  AND2_X1 U665 ( .A1(n573), .A2(n742), .ZN(n574) );
  OR2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U667 ( .A(KEYINPUT89), .ZN(n576) );
  XNOR2_X1 U668 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U669 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U670 ( .A1(n691), .A2(n608), .ZN(n582) );
  XNOR2_X1 U671 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n581) );
  XNOR2_X1 U672 ( .A(n582), .B(n581), .ZN(n585) );
  INV_X1 U673 ( .A(n583), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U675 ( .A(KEYINPUT35), .ZN(n586) );
  AND2_X1 U676 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U677 ( .A(KEYINPUT66), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(KEYINPUT22), .ZN(n592) );
  INV_X1 U679 ( .A(n676), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n595), .A2(n605), .ZN(n596) );
  NOR2_X1 U681 ( .A1(n670), .A2(n596), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n599), .A2(n597), .ZN(n632) );
  XNOR2_X1 U683 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n602), .A2(n642), .ZN(n604) );
  INV_X1 U685 ( .A(KEYINPUT94), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n678), .A2(n608), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n609) );
  NOR2_X1 U688 ( .A1(n611), .A2(n676), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT93), .ZN(n644) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT96), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT80), .B(n615), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n670), .A2(n595), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT104), .ZN(n759) );
  INV_X1 U695 ( .A(KEYINPUT45), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n729), .A2(G472), .ZN(n628) );
  XNOR2_X1 U697 ( .A(KEYINPUT84), .B(KEYINPUT62), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n628), .B(n363), .ZN(n630) );
  INV_X1 U699 ( .A(G952), .ZN(n629) );
  AND2_X1 U700 ( .A1(n629), .A2(G953), .ZN(n734) );
  NAND2_X1 U701 ( .A1(n630), .A2(n389), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n631), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U703 ( .A(n632), .B(G110), .ZN(G12) );
  XOR2_X1 U704 ( .A(G122), .B(KEYINPUT127), .Z(n634) );
  XNOR2_X1 U705 ( .A(n633), .B(n634), .ZN(G24) );
  NAND2_X1 U706 ( .A1(n729), .A2(G475), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT59), .B(KEYINPUT85), .Z(n635) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n639), .A2(n389), .ZN(n641) );
  XNOR2_X1 U710 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(G60) );
  XNOR2_X1 U712 ( .A(n642), .B(G119), .ZN(G21) );
  NAND2_X1 U713 ( .A1(n644), .A2(n656), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(G104), .ZN(G6) );
  XOR2_X1 U715 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U716 ( .A1(n644), .A2(n660), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(G107), .B(n647), .ZN(G9) );
  XOR2_X1 U719 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U720 ( .A1(n652), .A2(n660), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U722 ( .A(G128), .B(n650), .Z(G30) );
  XOR2_X1 U723 ( .A(G143), .B(n651), .Z(G45) );
  XOR2_X1 U724 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n654) );
  NAND2_X1 U725 ( .A1(n652), .A2(n656), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(G146), .B(n655), .ZN(G48) );
  NAND2_X1 U728 ( .A1(n659), .A2(n656), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT114), .ZN(n658) );
  XNOR2_X1 U730 ( .A(G113), .B(n658), .ZN(G15) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n661), .B(G116), .ZN(G18) );
  XNOR2_X1 U733 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U735 ( .A(G125), .B(n664), .ZN(G27) );
  XOR2_X1 U736 ( .A(G134), .B(n665), .Z(G36) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n668) );
  NAND2_X1 U738 ( .A1(n595), .A2(n666), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n669), .A2(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U746 ( .A(n679), .B(KEYINPUT51), .Z(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT118), .B(n680), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n699), .A2(n681), .ZN(n695) );
  NOR2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT119), .B(n686), .Z(n690) );
  NOR2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n693) );
  INV_X1 U754 ( .A(n691), .ZN(n692) );
  NOR2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n703) );
  INV_X1 U759 ( .A(n699), .ZN(n700) );
  NAND2_X1 U760 ( .A1(n700), .A2(n350), .ZN(n701) );
  NAND2_X1 U761 ( .A1(n701), .A2(n754), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n708) );
  INV_X1 U763 ( .A(n349), .ZN(n706) );
  INV_X1 U764 ( .A(KEYINPUT78), .ZN(n709) );
  INV_X1 U765 ( .A(KEYINPUT2), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n709), .A2(n704), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n712) );
  XNOR2_X1 U769 ( .A(n349), .B(n709), .ZN(n710) );
  NOR2_X1 U770 ( .A1(n710), .A2(KEYINPUT2), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U773 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n715) );
  XNOR2_X1 U774 ( .A(KEYINPUT79), .B(KEYINPUT55), .ZN(n714) );
  XNOR2_X1 U775 ( .A(n715), .B(n714), .ZN(n717) );
  XOR2_X1 U776 ( .A(n717), .B(n716), .Z(n718) );
  NAND2_X1 U777 ( .A1(n725), .A2(G469), .ZN(n723) );
  XOR2_X1 U778 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n720) );
  XNOR2_X1 U779 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n719) );
  XNOR2_X1 U780 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n734), .A2(n724), .ZN(G54) );
  NAND2_X1 U783 ( .A1(n725), .A2(G478), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n728), .A2(n734), .ZN(G63) );
  NAND2_X1 U786 ( .A1(n725), .A2(G217), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n734), .A2(n733), .ZN(G66) );
  OR2_X1 U788 ( .A1(n735), .A2(G953), .ZN(n739) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n740), .B(n741), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(G69) );
  XOR2_X1 U796 ( .A(n747), .B(n746), .Z(n751) );
  XOR2_X1 U797 ( .A(G227), .B(n751), .Z(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U799 ( .A1(G953), .A2(n749), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U801 ( .A(n751), .B(KEYINPUT125), .ZN(n753) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(G72) );
  XNOR2_X1 U805 ( .A(G140), .B(n758), .ZN(G42) );
  XNOR2_X1 U806 ( .A(G101), .B(n759), .ZN(G3) );
  XOR2_X1 U807 ( .A(n760), .B(G137), .Z(G39) );
  XOR2_X1 U808 ( .A(n761), .B(G131), .Z(G33) );
endmodule

