//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n461), .A2(G136), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n460), .A2(new_n462), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G162));
  OR2_X1    g052(.A1(new_n458), .A2(new_n459), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G126), .A3(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n462), .A2(KEYINPUT67), .A3(G138), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(KEYINPUT4), .C1(new_n459), .C2(new_n458), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n460), .B2(new_n480), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n479), .A2(new_n482), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G164));
  INV_X1    g063(.A(G62), .ZN(new_n489));
  INV_X1    g064(.A(G543), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .A3(G543), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n495), .B2(KEYINPUT69), .ZN(new_n498));
  OAI21_X1  g073(.A(G651), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n492), .A2(new_n494), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(G303));
  INV_X1    g080(.A(G303), .ZN(G166));
  NAND3_X1  g081(.A1(new_n500), .A2(G89), .A3(new_n502), .ZN(new_n507));
  NAND3_X1  g082(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT7), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n490), .B1(new_n502), .B2(KEYINPUT70), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n515), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n524), .A3(new_n515), .A4(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(G51), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n500), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n514), .A2(new_n527), .A3(new_n529), .ZN(G168));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(G52), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n520), .A2(new_n524), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT71), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n533), .B2(new_n525), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n492), .A2(new_n494), .B1(new_n517), .B2(new_n519), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G171));
  OAI21_X1  g115(.A(G43), .B1(new_n521), .B2(new_n526), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n492), .B2(new_n494), .ZN(new_n543));
  AND2_X1   g118(.A1(G68), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n547), .B(G651), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n535), .A2(G81), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n541), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n492), .B2(new_n494), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  INV_X1    g135(.A(G78), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n561), .B2(new_n490), .ZN(new_n562));
  NAND3_X1  g137(.A1(KEYINPUT75), .A2(G78), .A3(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT76), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n567), .B(G651), .C1(new_n559), .C2(new_n564), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n532), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n516), .A2(new_n572), .A3(G53), .A4(new_n520), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n535), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(G299));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n534), .B2(new_n539), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n534), .A2(KEYINPUT77), .A3(new_n539), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G301));
  NAND3_X1  g155(.A1(new_n514), .A2(new_n527), .A3(new_n529), .ZN(G286));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n492), .A2(new_n582), .A3(new_n494), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT80), .B1(new_n583), .B2(G651), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(KEYINPUT80), .A3(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n500), .A2(G87), .A3(new_n502), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n535), .A2(new_n589), .A3(G87), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n585), .A2(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n520), .A2(new_n524), .A3(G49), .A4(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n516), .A2(new_n594), .A3(G49), .A4(new_n520), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n535), .A2(G86), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n492), .B2(new_n494), .ZN(new_n602));
  AND2_X1   g177(.A1(G73), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g181(.A(KEYINPUT81), .B(G651), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G305));
  INV_X1    g184(.A(G47), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n533), .B2(new_n525), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n535), .A2(G85), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n538), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G290));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n500), .A2(new_n502), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n535), .A2(KEYINPUT10), .A3(G92), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n500), .A2(G66), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n620), .A2(new_n621), .B1(new_n624), .B2(G651), .ZN(new_n625));
  OAI21_X1  g200(.A(G54), .B1(new_n521), .B2(new_n526), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G301), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G284));
  AOI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G321));
  MUX2_X1   g206(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g207(.A(G299), .B(G286), .S(G868), .Z(G280));
  AND2_X1   g208(.A1(new_n625), .A2(new_n626), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT82), .B(G559), .Z(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(G860), .B2(new_n635), .ZN(G148));
  NOR2_X1   g211(.A1(new_n552), .A2(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT83), .Z(new_n639));
  AOI21_X1  g214(.A(new_n637), .B1(new_n639), .B2(G868), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n478), .A2(new_n463), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT13), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G2100), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT85), .Z(new_n647));
  AOI22_X1  g222(.A1(G123), .A2(new_n472), .B1(new_n461), .B2(G135), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n462), .A2(KEYINPUT86), .A3(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(KEYINPUT86), .B1(new_n462), .B2(G111), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n648), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  OAI211_X1 g228(.A(new_n647), .B(new_n653), .C1(G2100), .C2(new_n645), .ZN(G156));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT87), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n659), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(G14), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n666), .ZN(G401));
  XOR2_X1   g245(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT89), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n674), .B2(new_n671), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n680), .B(new_n682), .Z(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G32), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G105), .B2(new_n463), .ZN(new_n709));
  AOI22_X1  g284(.A1(G129), .A2(new_n472), .B1(new_n461), .B2(G141), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT27), .ZN(new_n714));
  INV_X1    g289(.A(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n461), .A2(G140), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n472), .A2(G128), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n462), .A2(G116), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n704), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n716), .A2(new_n728), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n730), .A2(KEYINPUT94), .A3(new_n462), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT94), .B1(new_n730), .B2(new_n462), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n733));
  NAND2_X1  g308(.A1(G103), .A2(G2104), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G2105), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n461), .A2(G139), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G33), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2072), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G35), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G162), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G2090), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(KEYINPUT101), .ZN(new_n746));
  NOR2_X1   g321(.A1(G4), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n634), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G1348), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n704), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n652), .B2(new_n704), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT98), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n704), .A2(G27), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT99), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n487), .B2(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n755), .A2(KEYINPUT98), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n757), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G34), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n765), .B2(G34), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n469), .A2(G29), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n762), .A2(new_n763), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n761), .B(new_n772), .C1(new_n744), .C2(G2090), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n729), .A2(new_n746), .A3(new_n750), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G16), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n775), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n745), .B2(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n775), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n775), .ZN(new_n782));
  AOI21_X1  g357(.A(KEYINPUT97), .B1(new_n782), .B2(G1966), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n777), .A2(new_n778), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(KEYINPUT97), .A3(G1966), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n775), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n552), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G16), .B2(G19), .ZN(new_n793));
  INV_X1    g368(.A(G1341), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n795), .B(new_n796), .C1(G1966), .C2(new_n782), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n774), .A2(new_n791), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n775), .A2(G23), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n593), .A2(new_n595), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n589), .B1(new_n535), .B2(G87), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n583), .A2(KEYINPUT80), .A3(G651), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n584), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(new_n775), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G6), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n608), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n775), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n775), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1971), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n814), .A2(KEYINPUT34), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n704), .A2(G25), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n461), .A2(G131), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n472), .A2(G119), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(new_n704), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT91), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G24), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n615), .B2(G16), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(G1986), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G1986), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n818), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n818), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT34), .B1(new_n814), .B2(new_n817), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n799), .B1(new_n841), .B2(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n798), .ZN(G150));
  NAND2_X1  g421(.A1(new_n634), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT102), .B(G55), .Z(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n521), .B2(new_n526), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n535), .A2(G93), .ZN(new_n851));
  AND2_X1   g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n500), .B2(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n853), .B2(new_n538), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n551), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n533), .A2(new_n525), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n858), .A2(G43), .B1(G81), .B2(new_n535), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n854), .B1(new_n858), .B2(new_n849), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n549), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n848), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n860), .A2(new_n866), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n711), .B(new_n721), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n487), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n738), .B2(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n875), .B2(new_n738), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n472), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n462), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G142), .B2(new_n461), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n644), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n825), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n889), .A3(new_n879), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n469), .B(new_n476), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n652), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g473(.A(new_n639), .B(new_n863), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(G299), .A2(new_n627), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n566), .A2(new_n568), .B1(G91), .B2(new_n535), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n903), .A2(new_n574), .B1(new_n625), .B2(new_n626), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(G299), .A2(new_n627), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(new_n574), .A3(new_n626), .A4(new_n625), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n902), .A2(new_n904), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n899), .ZN(new_n912));
  OAI22_X1  g487(.A1(new_n801), .A2(new_n805), .B1(new_n611), .B2(new_n614), .ZN(new_n913));
  OAI21_X1  g488(.A(G47), .B1(new_n521), .B2(new_n526), .ZN(new_n914));
  INV_X1    g489(.A(new_n614), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n591), .A2(new_n914), .A3(new_n915), .A4(new_n596), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT106), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(G305), .A2(G303), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n608), .A2(new_n504), .A3(new_n499), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G303), .B(new_n608), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n913), .A2(new_n916), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT107), .A3(KEYINPUT42), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n912), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n912), .B1(new_n933), .B2(new_n929), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n860), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n860), .ZN(G331));
  NAND2_X1  g513(.A1(new_n905), .A2(new_n909), .ZN(new_n939));
  INV_X1    g514(.A(new_n539), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT77), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n521), .A2(new_n526), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n531), .ZN(new_n943));
  AOI21_X1  g518(.A(G286), .B1(new_n577), .B2(new_n943), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n512), .A2(new_n513), .B1(new_n500), .B2(new_n528), .ZN(new_n945));
  AOI21_X1  g520(.A(G171), .B1(new_n527), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n857), .B(new_n861), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(G168), .B1(new_n578), .B2(new_n579), .ZN(new_n948));
  OAI21_X1  g523(.A(G286), .B1(new_n534), .B2(new_n539), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n862), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n939), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n906), .A2(new_n907), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n947), .B2(new_n950), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n927), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n911), .A2(new_n901), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n908), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n947), .A2(new_n956), .A3(new_n950), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n953), .B2(KEYINPUT109), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n960), .B(new_n952), .C1(new_n947), .C2(new_n950), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n928), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n948), .A2(new_n862), .A3(new_n949), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n862), .B1(new_n948), .B2(new_n949), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n911), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n939), .A2(new_n947), .A3(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n927), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G37), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n927), .B1(new_n972), .B2(KEYINPUT108), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT108), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT110), .B(new_n964), .C1(new_n975), .C2(new_n963), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n955), .A2(new_n962), .A3(new_n977), .A4(new_n963), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n955), .A2(new_n962), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT111), .B1(new_n981), .B2(new_n963), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n983), .A3(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n963), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(KEYINPUT44), .B2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n487), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n464), .A2(G40), .A3(new_n468), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n721), .B(new_n727), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n712), .A2(G1996), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n711), .A2(new_n715), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n824), .B(new_n827), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(G290), .A2(G1986), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n991), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n487), .A2(new_n988), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n487), .A2(new_n1005), .A3(new_n988), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1006), .A3(new_n990), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n1007), .A2(new_n1008), .A3(G2067), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n464), .A2(G40), .A3(new_n468), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n749), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1008), .B1(new_n1007), .B2(G2067), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT118), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1009), .A2(new_n1015), .A3(new_n1019), .A4(new_n1016), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n634), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  XNOR2_X1  g597(.A(G299), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n990), .B1(new_n1003), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n989), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT56), .B(G2072), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1006), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1005), .B1(new_n487), .B2(new_n988), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n990), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1956), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1024), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1021), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1038), .B(new_n1023), .C1(new_n1040), .C2(G1956), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1040), .B2(G1956), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT120), .B1(new_n1043), .B2(new_n1024), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1041), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT61), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1043), .A2(KEYINPUT120), .A3(new_n1024), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT121), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1046), .A2(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1048), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1007), .A2(new_n1008), .A3(G2067), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n749), .B2(new_n1014), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1019), .B1(new_n1055), .B2(new_n1016), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1020), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1051), .B(new_n1053), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1007), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1026), .A2(new_n989), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(G1996), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1027), .A2(new_n715), .B1(new_n1007), .B2(new_n1061), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n551), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1060), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1058), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1042), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1027), .A2(new_n757), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1014), .A2(new_n778), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1027), .A2(KEYINPUT53), .A3(new_n757), .ZN(new_n1077));
  AND4_X1   g652(.A1(G301), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1073), .A2(new_n1074), .B1(new_n1014), .B2(new_n778), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1026), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT123), .A3(new_n757), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT53), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT123), .B1(new_n1080), .B2(new_n757), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n629), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT125), .B1(new_n1085), .B2(KEYINPUT54), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1083), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n1081), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1090), .B2(new_n1079), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1087), .B(new_n1088), .C1(new_n1091), .C2(new_n1078), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1007), .A2(G8), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n608), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n604), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT115), .B(G86), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n599), .B1(new_n618), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(KEYINPUT49), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1094), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n806), .A2(G1976), .ZN(new_n1106));
  INV_X1    g681(.A(G1976), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(G288), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1094), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(G8), .A3(new_n1007), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1105), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G303), .A2(G8), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G2090), .ZN(new_n1116));
  INV_X1    g691(.A(G1971), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1040), .A2(new_n1116), .B1(new_n1063), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G8), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1115), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1014), .A2(G2090), .B1(new_n1027), .B2(G1971), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(G8), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1011), .A2(new_n769), .A3(new_n1013), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(G168), .C1(new_n1080), .C2(G1966), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1119), .A2(KEYINPUT122), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(KEYINPUT51), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT51), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1080), .A2(G1966), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1127), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1130), .A2(new_n1131), .B1(G168), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1088), .B1(new_n1136), .B2(G171), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n629), .B2(new_n1084), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1112), .A2(new_n1120), .A3(KEYINPUT126), .A4(new_n1123), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1126), .A2(new_n1135), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1072), .A2(new_n1093), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g718(.A(KEYINPUT62), .B1(G168), .B2(new_n1134), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1145), .A2(new_n1091), .A3(new_n1126), .A4(new_n1139), .ZN(new_n1146));
  OAI211_X1 g721(.A(G8), .B(G168), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(KEYINPUT63), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(new_n1112), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1105), .A2(new_n1107), .A3(new_n806), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1096), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1094), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1105), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1105), .A2(new_n1109), .A3(KEYINPUT116), .A4(new_n1111), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1149), .B(new_n1152), .C1(new_n1157), .C2(new_n1123), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1121), .B1(G8), .B2(new_n1122), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n1147), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1146), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1002), .B1(new_n1141), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n996), .A2(new_n998), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n991), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1001), .A2(KEYINPUT48), .A3(new_n991), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT48), .B1(new_n1001), .B2(new_n991), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n825), .A2(new_n827), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n995), .A2(new_n1173), .B1(G2067), .B2(new_n721), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n991), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n991), .A2(new_n715), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1177));
  INV_X1    g752(.A(new_n992), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n991), .B1(new_n1178), .B2(new_n711), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT127), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1175), .B1(new_n1181), .B2(KEYINPUT47), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1172), .B(new_n1182), .C1(KEYINPUT47), .C2(new_n1181), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(G319), .ZN(new_n1186));
  NOR3_X1   g760(.A1(G401), .A2(new_n1186), .A3(G227), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n702), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n894), .B2(new_n896), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n1189), .A2(new_n976), .A3(new_n978), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


