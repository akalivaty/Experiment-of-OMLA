//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT66), .B(G131), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT70), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G237), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G214), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(G237), .B1(new_n191), .B2(new_n193), .ZN(new_n199));
  AOI21_X1  g013(.A(G143), .B1(new_n199), .B2(G214), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n189), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n187), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n197), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n188), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n202), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n210), .B1(new_n214), .B2(new_n208), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(G146), .B(new_n210), .C1(new_n214), .C2(new_n208), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n204), .A2(new_n205), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(KEYINPUT89), .A3(KEYINPUT17), .A4(new_n189), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n203), .A2(new_n207), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n204), .A2(KEYINPUT18), .A3(G131), .A4(new_n205), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(G146), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n213), .A3(new_n216), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G113), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n223), .A2(new_n236), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G475), .ZN(new_n243));
  NOR2_X1   g057(.A1(G475), .A2(G902), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n226), .A2(new_n227), .B1(new_n230), .B2(new_n229), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n214), .B(KEYINPUT19), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n218), .B1(new_n250), .B2(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n201), .B2(new_n206), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n237), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n239), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n244), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n239), .B2(new_n253), .ZN(new_n256));
  OAI22_X1  g070(.A1(KEYINPUT91), .A2(new_n254), .B1(new_n256), .B2(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n243), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT92), .ZN(new_n262));
  INV_X1    g076(.A(G122), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT92), .A2(G122), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(G116), .ZN(new_n267));
  OR3_X1    g081(.A1(new_n266), .A2(KEYINPUT93), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n265), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT92), .A2(G122), .ZN(new_n270));
  OAI21_X1  g084(.A(G116), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n267), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT93), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n274), .A3(G107), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n197), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT13), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT94), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT94), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n197), .A2(KEYINPUT13), .A3(G128), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n281), .A4(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n283), .B1(new_n290), .B2(G134), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n277), .A2(new_n278), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n282), .B1(new_n279), .B2(new_n281), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT14), .ZN(new_n295));
  OAI21_X1  g109(.A(G107), .B1(new_n266), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n273), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n271), .A2(new_n295), .A3(G107), .A4(new_n272), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI211_X1 g115(.A(KEYINPUT95), .B(new_n294), .C1(new_n297), .C2(new_n298), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT9), .B(G234), .Z(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(G217), .A3(new_n190), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n307));
  INV_X1    g121(.A(new_n305), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n292), .B(new_n308), .C1(new_n301), .C2(new_n302), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n303), .A2(KEYINPUT96), .A3(new_n305), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n241), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G478), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT15), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G952), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G953), .ZN(new_n317));
  INV_X1    g131(.A(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n195), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n241), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n314), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n310), .A2(new_n241), .A3(new_n311), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n315), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n260), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G217), .B1(new_n318), .B2(G902), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT73), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G128), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT68), .B(G119), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(new_n280), .ZN(new_n335));
  OR2_X1    g149(.A1(KEYINPUT24), .A2(G110), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT24), .A2(G110), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(KEYINPUT24), .A2(G110), .ZN(new_n340));
  NOR2_X1   g154(.A1(KEYINPUT24), .A2(G110), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT74), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n330), .B1(new_n335), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n331), .A2(KEYINPUT68), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n332), .B1(new_n348), .B2(G128), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n339), .A4(new_n342), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT23), .B(new_n333), .C1(new_n334), .C2(new_n280), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n334), .A2(new_n353), .A3(new_n280), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(G110), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n219), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G110), .B1(new_n352), .B2(new_n354), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n335), .A2(new_n343), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n218), .B(new_n230), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n356), .B2(new_n359), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(new_n365), .B2(new_n241), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  NOR4_X1   g181(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(G902), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n329), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT76), .B(new_n329), .C1(new_n366), .C2(new_n368), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n329), .A2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n327), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n235), .A2(KEYINPUT79), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n276), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(G104), .B2(G107), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT3), .A2(G107), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n235), .A2(KEYINPUT79), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n276), .A3(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT3), .A2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT80), .B1(new_n396), .B2(new_n385), .ZN(new_n397));
  INV_X1    g211(.A(new_n388), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n382), .B2(new_n383), .ZN(new_n399));
  AND2_X1   g213(.A1(KEYINPUT3), .A2(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(G104), .B2(new_n388), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n399), .A2(KEYINPUT80), .A3(new_n401), .A4(new_n385), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n387), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(KEYINPUT2), .A2(G113), .ZN(new_n405));
  NOR2_X1   g219(.A1(KEYINPUT2), .A2(G113), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n261), .A2(G119), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n407), .B(new_n408), .C1(new_n334), .C2(new_n261), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n348), .A2(G116), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(KEYINPUT69), .A3(new_n408), .A4(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n346), .A2(G119), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n331), .A2(KEYINPUT68), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(G116), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT5), .B(new_n408), .C1(new_n334), .C2(new_n261), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n348), .A2(KEYINPUT84), .A3(new_n415), .A4(G116), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n420), .A2(G113), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n404), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n399), .A2(new_n385), .A3(new_n401), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n402), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(new_n387), .A3(new_n414), .A4(new_n423), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n429), .A2(new_n402), .B1(new_n384), .B2(new_n386), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT86), .A3(new_n414), .A4(new_n423), .ZN(new_n434));
  XOR2_X1   g248(.A(G110), .B(G122), .Z(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT8), .Z(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n216), .A2(G143), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n197), .A2(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT0), .A2(G128), .ZN(new_n441));
  OR2_X1    g255(.A1(KEYINPUT0), .A2(G128), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n216), .A3(G143), .ZN(new_n445));
  INV_X1    g259(.A(new_n441), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT64), .B1(new_n197), .B2(G146), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n197), .A2(G146), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT65), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n444), .B1(new_n216), .B2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n438), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n445), .A4(new_n446), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n443), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(new_n212), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n445), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT1), .ZN(new_n459));
  OAI21_X1  g273(.A(G128), .B1(new_n448), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n440), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n461), .A3(new_n212), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n190), .A2(G224), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n456), .A2(new_n462), .B1(KEYINPUT7), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n462), .C1(new_n455), .C2(new_n212), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n437), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n437), .A2(new_n468), .A3(KEYINPUT87), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n412), .A2(new_n408), .ZN(new_n473));
  INV_X1    g287(.A(new_n407), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n411), .A2(new_n413), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n399), .A2(new_n401), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n429), .A2(new_n402), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT81), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n477), .A2(new_n480), .A3(KEYINPUT4), .A4(G101), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(G101), .C1(new_n391), .C2(new_n395), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n476), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n435), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n431), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n471), .A2(new_n472), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n456), .A2(new_n462), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(new_n463), .Z(new_n491));
  XNOR2_X1  g305(.A(new_n482), .B(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n429), .A2(new_n402), .A3(new_n478), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n475), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n404), .A2(new_n424), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n435), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n488), .A3(KEYINPUT6), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n487), .B1(new_n486), .B2(new_n431), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT85), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n499), .B(new_n435), .C1(new_n494), .C2(new_n495), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n491), .B(new_n497), .C1(new_n500), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n489), .A2(new_n241), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n507), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n489), .A2(new_n504), .A3(new_n241), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n380), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n304), .ZN(new_n512));
  OAI21_X1  g326(.A(G221), .B1(new_n512), .B2(G902), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT77), .ZN(new_n514));
  INV_X1    g328(.A(G469), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT11), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n282), .B2(G137), .ZN(new_n517));
  INV_X1    g331(.A(G137), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT11), .A3(G134), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n282), .A2(G137), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G131), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n188), .A2(new_n517), .A3(new_n519), .A4(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT82), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n458), .A2(new_n461), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n433), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n452), .A2(new_n445), .ZN(new_n529));
  INV_X1    g343(.A(new_n460), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n458), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n387), .C1(new_n397), .C2(new_n403), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n526), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT12), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n455), .B1(new_n479), .B2(new_n485), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n433), .A2(KEYINPUT10), .A3(new_n527), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(new_n538), .A3(new_n525), .A4(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(G110), .B(G140), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT78), .ZN(new_n542));
  INV_X1    g356(.A(new_n194), .ZN(new_n543));
  INV_X1    g357(.A(G227), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n542), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n526), .C1(new_n528), .C2(new_n533), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n535), .A2(new_n540), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n551), .B2(new_n540), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n549), .B1(new_n552), .B2(KEYINPUT83), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n554), .B(new_n546), .C1(new_n551), .C2(new_n540), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n515), .B(new_n241), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n515), .A2(new_n241), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n535), .A2(new_n540), .A3(new_n548), .ZN(new_n558));
  INV_X1    g372(.A(new_n546), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n540), .A2(new_n546), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n557), .B1(new_n561), .B2(G469), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n514), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n450), .A2(new_n454), .ZN(new_n564));
  INV_X1    g378(.A(new_n443), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n524), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n518), .A2(G134), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n225), .B1(new_n567), .B2(new_n520), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT67), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n527), .A2(new_n523), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n475), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n566), .A2(new_n572), .A3(KEYINPUT30), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT30), .B1(new_n566), .B2(new_n572), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n577), .B2(new_n476), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n199), .A2(G210), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT28), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n566), .A2(new_n572), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n476), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n589), .B2(new_n573), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n573), .A2(new_n587), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n586), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT30), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n566), .A2(new_n572), .A3(KEYINPUT30), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n476), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n579), .A3(new_n573), .A4(new_n584), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT31), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n585), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(G472), .A2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT32), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n597), .A2(new_n573), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n586), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT29), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n475), .B1(new_n566), .B2(new_n572), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT28), .B1(new_n574), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n591), .A3(new_n584), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n241), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT72), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n609), .B2(new_n591), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n590), .A2(KEYINPUT72), .ZN(new_n615));
  NOR4_X1   g429(.A1(new_n614), .A2(new_n615), .A3(new_n607), .A4(new_n586), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n600), .A2(KEYINPUT32), .A3(new_n601), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n604), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n378), .A2(new_n511), .A3(new_n563), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NAND2_X1  g435(.A1(new_n501), .A2(new_n502), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n498), .A2(KEYINPUT85), .A3(new_n499), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n498), .A2(new_n499), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(new_n488), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n491), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n509), .B1(new_n626), .B2(new_n489), .ZN(new_n627));
  INV_X1    g441(.A(new_n510), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n379), .B(new_n323), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n303), .A2(new_n631), .A3(new_n305), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n303), .B2(new_n305), .ZN(new_n633));
  OAI211_X1 g447(.A(KEYINPUT33), .B(new_n309), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n310), .A2(new_n635), .A3(new_n311), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n313), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n312), .A2(new_n313), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n260), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n630), .A2(KEYINPUT98), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n629), .B2(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n600), .A2(new_n241), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n646), .A2(G472), .B1(new_n600), .B2(new_n601), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n563), .A2(new_n376), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND2_X1  g466(.A1(new_n315), .A2(new_n325), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n239), .A2(new_n253), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n244), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT20), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n256), .A2(new_n246), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n242), .A2(KEYINPUT99), .A3(G475), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  AOI21_X1  g474(.A(G902), .B1(new_n238), .B2(new_n239), .ZN(new_n661));
  INV_X1    g475(.A(G475), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n649), .A2(new_n630), .A3(new_n653), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G107), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n508), .A2(new_n510), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n563), .A2(new_n669), .A3(new_n379), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n356), .A2(new_n359), .ZN(new_n671));
  INV_X1    g485(.A(new_n362), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT36), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n373), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n371), .A2(new_n372), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n371), .A2(new_n681), .A3(new_n678), .A4(new_n372), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n680), .A2(new_n327), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n670), .A2(new_n647), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n682), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n319), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n320), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n658), .A2(new_n659), .A3(new_n663), .A4(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n325), .B2(new_n315), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n670), .A2(new_n619), .A3(new_n688), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XNOR2_X1  g510(.A(new_n691), .B(KEYINPUT39), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n563), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n627), .A2(new_n628), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n703), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n669), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n604), .A2(new_n618), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n578), .A2(new_n586), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n574), .A2(new_n608), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n710), .B2(new_n586), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n260), .A2(new_n379), .A3(new_n653), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n688), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n701), .A2(new_n707), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT105), .B(G143), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G45));
  AND3_X1   g533(.A1(new_n260), .A2(new_n640), .A3(new_n692), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n670), .A2(new_n619), .A3(new_n688), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  AND2_X1   g536(.A1(new_n619), .A2(new_n376), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n241), .B1(new_n553), .B2(new_n555), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n515), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI221_X1 g541(.A(new_n241), .B1(new_n725), .B2(new_n515), .C1(new_n553), .C2(new_n555), .ZN(new_n728));
  INV_X1    g542(.A(new_n514), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n643), .A2(new_n645), .A3(new_n723), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND3_X1  g548(.A1(new_n376), .A2(new_n664), .A3(new_n653), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n629), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n379), .B1(new_n627), .B2(new_n628), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n730), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n619), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n619), .A3(new_n683), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NOR2_X1   g556(.A1(new_n702), .A2(new_n715), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n586), .B1(new_n614), .B2(new_n615), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n599), .A3(new_n585), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n646), .A2(G472), .B1(new_n745), .B2(new_n601), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n376), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n731), .A3(new_n748), .A4(new_n323), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT107), .B(G122), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G24));
  AND3_X1   g565(.A1(new_n680), .A2(new_n746), .A3(new_n682), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n738), .A2(new_n720), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NAND2_X1  g568(.A1(new_n556), .A2(new_n562), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n729), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n508), .A2(new_n379), .A3(new_n510), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n723), .A3(new_n720), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n619), .A2(new_n376), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n756), .A3(new_n757), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT42), .A3(new_n720), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  AND3_X1   g580(.A1(new_n758), .A2(new_n723), .A3(new_n694), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT108), .B(G134), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G36));
  INV_X1    g583(.A(new_n260), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n640), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT43), .A3(new_n640), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n647), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n688), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n757), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n776), .A4(new_n688), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n561), .A2(KEYINPUT45), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(G469), .B1(new_n561), .B2(KEYINPUT45), .ZN(new_n783));
  OAI22_X1  g597(.A1(new_n782), .A2(new_n783), .B1(new_n515), .B2(new_n241), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n556), .B1(new_n784), .B2(new_n785), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n729), .B(new_n698), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n779), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  XNOR2_X1  g606(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n729), .B(new_n793), .C1(new_n787), .C2(new_n788), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n720), .A2(new_n375), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n619), .A3(new_n757), .ZN(new_n796));
  INV_X1    g610(.A(new_n788), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n514), .B1(new_n797), .B2(new_n786), .ZN(new_n798));
  NOR2_X1   g612(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n794), .B(new_n796), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR2_X1   g615(.A1(new_n707), .A2(new_n714), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n376), .A2(new_n379), .A3(new_n729), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n727), .A2(new_n728), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n771), .B(new_n803), .C1(KEYINPUT49), .C2(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n802), .B(new_n805), .C1(KEYINPUT49), .C2(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n511), .A2(new_n563), .A3(new_n619), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n511), .A2(new_n563), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n680), .A2(new_n327), .A3(new_n647), .A4(new_n682), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n807), .A2(new_n377), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n656), .A3(new_n258), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n653), .A2(new_n812), .A3(new_n243), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n641), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n648), .A2(new_n814), .A3(new_n629), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n619), .B(new_n738), .C1(new_n736), .C2(new_n683), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n732), .A3(new_n749), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n767), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n720), .A2(new_n680), .A3(new_n682), .A4(new_n746), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n693), .A2(new_n653), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n619), .A3(new_n680), .A4(new_n682), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n758), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT42), .B1(new_n763), .B2(new_n720), .ZN(new_n825));
  AND4_X1   g639(.A1(KEYINPUT42), .A2(new_n758), .A3(new_n720), .A4(new_n723), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n819), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n807), .A2(new_n687), .ZN(new_n829));
  INV_X1    g643(.A(new_n820), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n829), .A2(new_n694), .B1(new_n830), .B2(new_n738), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n679), .A2(new_n691), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n743), .A2(new_n714), .A3(new_n563), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n721), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n695), .A2(new_n721), .A3(new_n753), .A4(new_n833), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n739), .A2(new_n741), .A3(new_n749), .ZN(new_n840));
  INV_X1    g654(.A(new_n814), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n649), .A2(new_n630), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n684), .A3(new_n620), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n767), .B1(new_n761), .B2(new_n764), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n732), .A4(new_n824), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n834), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n835), .A2(KEYINPUT110), .A3(new_n836), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n839), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n835), .A2(new_n836), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n847), .B2(new_n837), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT53), .B(new_n828), .C1(new_n858), .C2(new_n850), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n828), .A2(new_n838), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g677(.A(KEYINPUT111), .B(KEYINPUT53), .C1(new_n828), .C2(new_n838), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n856), .B(new_n859), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n380), .B1(KEYINPUT114), .B2(KEYINPUT50), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n704), .A2(new_n706), .A3(new_n730), .A4(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n775), .A2(KEYINPUT113), .A3(new_n689), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT113), .B1(new_n775), .B2(new_n689), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n748), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n870), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n775), .A2(KEYINPUT113), .A3(new_n689), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n747), .B(new_n757), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n798), .A2(new_n799), .ZN(new_n877));
  INV_X1    g691(.A(new_n794), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n877), .A2(new_n878), .B1(new_n729), .B2(new_n804), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n714), .A2(new_n375), .A3(new_n319), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n730), .A2(new_n757), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT115), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n260), .A2(new_n640), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n752), .B(new_n882), .C1(new_n869), .C2(new_n870), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n873), .A2(new_n880), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n895));
  OAI221_X1 g709(.A(new_n895), .B1(new_n729), .B2(new_n804), .C1(new_n877), .C2(new_n878), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n876), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n873), .A4(new_n890), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n738), .B(new_n748), .C1(new_n869), .C2(new_n870), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n884), .A2(new_n642), .A3(new_n886), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n317), .A4(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n723), .B(new_n882), .C1(new_n869), .C2(new_n870), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT48), .Z(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n893), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT118), .B1(new_n866), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n854), .A3(KEYINPUT118), .A4(new_n865), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n316), .A2(new_n190), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n806), .B1(new_n909), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n194), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G902), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n509), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n625), .B(new_n491), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n915), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n834), .A2(new_n837), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n862), .B1(new_n924), .B2(new_n846), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT111), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n861), .A2(new_n860), .A3(new_n862), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n241), .B1(new_n928), .B2(new_n859), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n507), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n930), .B2(new_n916), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n923), .A2(new_n931), .ZN(G51));
  XNOR2_X1  g746(.A(new_n557), .B(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n856), .B1(new_n928), .B2(new_n859), .ZN(new_n934));
  INV_X1    g748(.A(new_n865), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n553), .A2(new_n555), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g752(.A1(new_n918), .A2(new_n782), .A3(new_n783), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n914), .B1(new_n938), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n239), .B(new_n253), .C1(new_n918), .C2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(new_n654), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n915), .ZN(G60));
  NAND2_X1  g758(.A1(new_n634), .A2(new_n636), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT119), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n854), .A2(new_n865), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT59), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n917), .A2(new_n855), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n865), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n950), .A2(new_n914), .A3(new_n953), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n917), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n671), .A2(new_n672), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n917), .A2(new_n674), .A3(new_n675), .A4(new_n958), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n915), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n915), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  AOI21_X1  g783(.A(new_n190), .B1(new_n322), .B2(G224), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT122), .Z(new_n971));
  INV_X1    g785(.A(new_n818), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n543), .ZN(new_n973));
  INV_X1    g787(.A(new_n625), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(G898), .B2(new_n194), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  OAI21_X1  g790(.A(new_n543), .B1(new_n544), .B2(new_n690), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT126), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n577), .B(new_n250), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n194), .A2(G900), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n695), .A2(new_n721), .A3(new_n753), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n791), .A2(new_n800), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n790), .A2(new_n723), .A3(new_n743), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n986), .A2(new_n987), .A3(new_n845), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n983), .B1(new_n989), .B2(new_n194), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n984), .A2(KEYINPUT123), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n984), .A2(KEYINPUT123), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n791), .A2(new_n988), .A3(new_n800), .A4(new_n845), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(new_n543), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT124), .B1(new_n998), .B2(new_n983), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n992), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n986), .A2(new_n717), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n986), .A2(KEYINPUT62), .A3(new_n717), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OR4_X1    g819(.A1(new_n699), .A2(new_n814), .A3(new_n762), .A4(new_n757), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n987), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n982), .A2(new_n194), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n979), .B(new_n981), .C1(new_n1000), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n981), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n992), .A2(new_n999), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n978), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  INV_X1    g831(.A(new_n606), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n605), .A2(new_n586), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n853), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1017), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n997), .B2(new_n972), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n578), .A2(new_n586), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n915), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1017), .B1(new_n1008), .B2(new_n818), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n1022), .B(new_n1026), .C1(new_n1027), .C2(new_n709), .ZN(G57));
endmodule


