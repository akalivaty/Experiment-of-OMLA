//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT67), .Z(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n462), .B2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n461), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(G126), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT3), .B(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n462), .B2(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT68), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n461), .B2(G114), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n485), .A2(new_n491), .A3(new_n494), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n512), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n514), .C2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n522), .A2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  XNOR2_X1  g104(.A(KEYINPUT72), .B(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n512), .A2(new_n530), .B1(new_n514), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n518), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n512), .A2(new_n536), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n518), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT73), .Z(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  AND2_X1   g122(.A1(new_n511), .A2(G65), .ZN(new_n548));
  AND2_X1   g123(.A1(G78), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(G53), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT74), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n521), .A2(G91), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n550), .A2(new_n556), .A3(new_n557), .ZN(G299));
  OR2_X1    g133(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  INV_X1    g135(.A(new_n514), .ZN(new_n561));
  AOI22_X1  g136(.A1(G87), .A2(new_n521), .B1(new_n561), .B2(G49), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(G288));
  NAND3_X1  g139(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n509), .B2(new_n510), .ZN(new_n569));
  AND2_X1   g144(.A1(G73), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  INV_X1    g149(.A(new_n511), .ZN(new_n575));
  INV_X1    g150(.A(G60), .ZN(new_n576));
  INV_X1    g151(.A(G72), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n508), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  OAI221_X1 g155(.A(new_n580), .B1(new_n577), .B2(new_n508), .C1(new_n575), .C2(new_n576), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(G651), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(G85), .A2(new_n521), .B1(new_n561), .B2(G47), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n582), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n506), .A2(G92), .A3(new_n511), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n575), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n561), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G286), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(G299), .B(KEYINPUT77), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G297));
  AOI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n541), .ZN(G323));
  XOR2_X1   g186(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n612));
  XNOR2_X1  g187(.A(G323), .B(new_n612), .ZN(G282));
  NAND2_X1  g188(.A1(new_n490), .A2(new_n468), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n473), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n475), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n461), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n618), .A2(new_n619), .A3(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n644), .B2(new_n646), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n651), .A2(new_n647), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n648), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n659), .A2(new_n664), .A3(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n663), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT83), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n671), .B(new_n675), .Z(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NOR2_X1   g252(.A1(G171), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G5), .B2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G1961), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT31), .B(G11), .Z(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(G28), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(G28), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G168), .A2(new_n677), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n677), .B2(G21), .ZN(new_n691));
  INV_X1    g266(.A(G1966), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n689), .B1(new_n683), .B2(new_n624), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n681), .B(new_n693), .C1(new_n692), .C2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT92), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n683), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n683), .ZN(new_n697));
  INV_X1    g272(.A(G2090), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G4), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n597), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1348), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n683), .A2(G26), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT88), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n708));
  INV_X1    g283(.A(G116), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n475), .B2(G140), .ZN(new_n711));
  AOI21_X1  g286(.A(KEYINPUT87), .B1(new_n473), .B2(G128), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n490), .A2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n714));
  INV_X1    g289(.A(G128), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n711), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n707), .B1(new_n717), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2067), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  INV_X1    g297(.A(G129), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n713), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n468), .A2(G105), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n461), .ZN(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(new_n683), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n683), .B2(G32), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G34), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G29), .B2(G160), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n731), .A2(new_n732), .B1(G2084), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n731), .A2(new_n732), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(G2084), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n704), .A2(new_n720), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n683), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n475), .A2(G139), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n472), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2105), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT89), .Z(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n742), .B1(new_n754), .B2(new_n683), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n683), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n683), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT93), .B(G2078), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n679), .A2(new_n680), .ZN(new_n762));
  INV_X1    g337(.A(G1341), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n541), .A2(new_n677), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n677), .B2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n761), .B(new_n766), .C1(new_n763), .C2(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n701), .A2(new_n741), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n677), .A2(G20), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT23), .Z(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n695), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n677), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(G288), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n677), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT85), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n677), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n677), .ZN(new_n783));
  INV_X1    g358(.A(G1971), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G6), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n573), .B2(G16), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n780), .A2(new_n781), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n677), .A2(G24), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT84), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G290), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1986), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT36), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n473), .A2(G119), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n475), .A2(G131), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n461), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n806));
  OR4_X1    g381(.A1(KEYINPUT86), .A2(new_n796), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT86), .B(KEYINPUT36), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n796), .B2(new_n806), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n774), .A2(new_n807), .A3(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n597), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  INV_X1    g388(.A(new_n541), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n521), .A2(G93), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n561), .A2(G55), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n815), .B(new_n816), .C1(new_n518), .C2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n813), .B(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n824), .A2(new_n825), .A3(G860), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n818), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(new_n802), .B(new_n615), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n729), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n717), .A2(G164), .ZN(new_n833));
  INV_X1    g408(.A(G140), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n461), .A2(G116), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n726), .A2(new_n834), .B1(new_n835), .B2(new_n708), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n473), .A2(KEYINPUT87), .A3(G128), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n502), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n832), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n717), .A2(G164), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n502), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n729), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n754), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n842), .A2(new_n843), .A3(new_n729), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n729), .B1(new_n842), .B2(new_n843), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT96), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n841), .B2(new_n844), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n752), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT96), .B1(new_n847), .B2(new_n848), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n841), .A2(new_n850), .A3(new_n844), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n855), .A2(new_n856), .B1(new_n751), .B2(new_n747), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n475), .A2(G142), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT98), .Z(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  INV_X1    g436(.A(G118), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(G2105), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n473), .B2(G130), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n854), .A2(new_n858), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n857), .A2(KEYINPUT97), .B1(new_n754), .B2(new_n845), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n852), .A2(new_n853), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n831), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n624), .B(G160), .Z(new_n872));
  XNOR2_X1  g447(.A(G162), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n865), .B1(new_n854), .B2(new_n858), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n869), .A3(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n830), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n871), .A2(KEYINPUT99), .A3(new_n873), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n873), .B1(new_n871), .B2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(G37), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n881), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(G395));
  NAND2_X1  g461(.A1(new_n818), .A2(new_n600), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G288), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n821), .B(new_n607), .ZN(new_n892));
  INV_X1    g467(.A(G299), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n596), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n596), .A2(new_n893), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT101), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT102), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n892), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n895), .B2(new_n897), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n903), .B1(new_n892), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n891), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n887), .B1(new_n910), .B2(new_n600), .ZN(G295));
  OAI21_X1  g486(.A(new_n887), .B1(new_n910), .B2(new_n600), .ZN(G331));
  NAND2_X1  g487(.A1(G301), .A2(KEYINPUT103), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g489(.A1(G168), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G286), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n822), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(G168), .B1(new_n913), .B2(new_n914), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n821), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n822), .A2(KEYINPUT104), .A3(new_n915), .A4(new_n917), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n895), .A2(new_n897), .A3(new_n905), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n925), .B(new_n928), .C1(new_n907), .C2(new_n927), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n921), .B(new_n918), .C1(new_n900), .C2(new_n902), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n890), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n918), .A2(new_n921), .ZN(new_n933));
  INV_X1    g508(.A(new_n906), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n926), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n923), .A2(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n899), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n890), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n931), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n907), .A2(new_n933), .B1(new_n936), .B2(new_n899), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n890), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n939), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n931), .A2(new_n940), .A3(KEYINPUT43), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n950), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n483), .A2(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT69), .B1(new_n497), .B2(G2105), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n495), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n956), .A2(new_n498), .B1(new_n493), .B2(KEYINPUT68), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n958), .B2(KEYINPUT45), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  AND4_X1   g535(.A1(new_n953), .A2(new_n502), .A3(KEYINPUT45), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n485), .A2(new_n491), .ZN(new_n963));
  NAND2_X1  g538(.A1(G126), .A2(G2105), .ZN(new_n964));
  OR2_X1    g539(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n965));
  NAND2_X1  g540(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n501), .B1(new_n967), .B2(new_n487), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n960), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n467), .A2(new_n469), .ZN(new_n972));
  INV_X1    g547(.A(G125), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n965), .B2(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(new_n465), .ZN(new_n975));
  OAI21_X1  g550(.A(G2105), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n976), .A3(G40), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT106), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n979));
  NAND3_X1  g554(.A1(G160), .A2(new_n979), .A3(G40), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n971), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n692), .B1(new_n962), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n502), .B2(new_n960), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n502), .A2(new_n984), .A3(new_n960), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2084), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n952), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G168), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT63), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n521), .A2(G86), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT110), .B(G1981), .Z(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n993), .A2(new_n571), .A3(new_n565), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n573), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n978), .A2(new_n980), .A3(new_n958), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n996), .B(KEYINPUT49), .C1(new_n573), .C2(new_n997), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1000), .A2(G8), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n776), .A2(G1976), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n1006), .A3(G8), .A4(new_n1001), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1001), .A2(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G288), .A2(new_n1005), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n991), .A2(new_n992), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n979), .B1(G160), .B2(G40), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n979), .A2(new_n972), .A3(new_n976), .A4(G40), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n971), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n784), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n502), .A2(new_n984), .A3(new_n960), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n978), .A3(new_n980), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1022), .B2(G2090), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n986), .A2(new_n985), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(KEYINPUT108), .A3(new_n1015), .A4(new_n698), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1012), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1028), .B(new_n1029), .Z(new_n1035));
  AOI22_X1  g610(.A1(new_n698), .A2(new_n987), .B1(new_n1017), .B2(new_n784), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n952), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1011), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1026), .A2(new_n1030), .A3(G8), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n992), .B1(new_n1040), .B2(new_n991), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(G1976), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1003), .A2(new_n1042), .B1(new_n573), .B2(new_n995), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1039), .A2(new_n1011), .B1(new_n1043), .B2(new_n1008), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT111), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n1046));
  OAI221_X1 g621(.A(new_n1046), .B1(new_n1043), .B2(new_n1008), .C1(new_n1039), .C2(new_n1011), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1034), .A2(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G286), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT118), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n982), .B2(new_n989), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n990), .A2(KEYINPUT51), .A3(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n990), .B2(KEYINPUT119), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n502), .B2(new_n960), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n983), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1016), .A2(KEYINPUT112), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n958), .A2(new_n953), .A3(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1966), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1022), .A2(G2084), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT119), .B(G8), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1053), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1050), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(new_n1062), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT120), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1052), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1956), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1022), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(new_n756), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1015), .A2(new_n971), .A3(new_n1016), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT114), .B1(new_n554), .B2(new_n555), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(KEYINPUT57), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G299), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n554), .A2(new_n555), .B1(new_n521), .B2(G91), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n550), .C1(new_n1079), .C2(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1348), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1022), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1001), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n719), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n596), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1084), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1075), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1091), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT117), .B(new_n1093), .C1(new_n1094), .C2(new_n1091), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1087), .A2(new_n1089), .A3(new_n596), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1084), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .A3(new_n1085), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1015), .A2(new_n1106), .A3(new_n971), .A4(new_n1016), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1001), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n814), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1086), .A2(new_n1022), .B1(new_n1088), .B2(new_n719), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n596), .A2(KEYINPUT60), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1110), .A2(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1101), .A2(new_n1105), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1092), .B1(new_n1099), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT124), .B(G2078), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1055), .B2(new_n977), .ZN(new_n1123));
  INV_X1    g698(.A(new_n977), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(KEYINPUT123), .C1(new_n958), .C2(KEYINPUT45), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1128), .B(new_n1121), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G2078), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1015), .A2(new_n1131), .A3(new_n971), .A4(new_n1016), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1133));
  AOI22_X1  g708(.A1(new_n1132), .A2(new_n1133), .B1(new_n680), .B2(new_n1022), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1130), .A2(new_n1135), .A3(G171), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1056), .A2(new_n1131), .A3(new_n1059), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT121), .A4(new_n1131), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT53), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1141), .B2(new_n1134), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1119), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1134), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1134), .B(KEYINPUT126), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(G171), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1135), .A2(G171), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1119), .B1(new_n1149), .B2(new_n1141), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1040), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1118), .A2(new_n1143), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1048), .B1(new_n1073), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT127), .B(new_n1048), .C1(new_n1073), .C2(new_n1152), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1052), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1053), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1071), .B2(KEYINPUT120), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT62), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1157), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1142), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1040), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1155), .A2(new_n1156), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n983), .A2(new_n971), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n729), .B(G1996), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n839), .B(G2067), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n802), .B(new_n804), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1170), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n1178), .A2(KEYINPUT107), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1170), .B1(new_n1178), .B2(KEYINPUT107), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1168), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1170), .B1(new_n729), .B2(new_n1172), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1170), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT46), .B1(new_n1170), .B2(G1996), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT47), .Z(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT48), .B1(new_n1179), .B2(new_n1169), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1176), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1179), .A2(KEYINPUT48), .A3(new_n1169), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n804), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n802), .A2(new_n1193), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n1173), .A2(new_n1194), .B1(G2067), .B2(new_n717), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1169), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1188), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1183), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g774(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1201));
  OAI21_X1  g775(.A(new_n1201), .B1(new_n948), .B2(new_n949), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n881), .B2(new_n883), .ZN(G308));
  NAND2_X1  g777(.A1(new_n881), .A2(new_n883), .ZN(new_n1204));
  OAI211_X1 g778(.A(new_n1204), .B(new_n1201), .C1(new_n949), .C2(new_n948), .ZN(G225));
endmodule


