//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(G43gat), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT92), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n217), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n209), .B1(new_n206), .B2(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT93), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(G29gat), .A3(G36gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n220), .A2(new_n205), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n219), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT94), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n219), .A3(KEYINPUT94), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n216), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n221), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n205), .A3(new_n220), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT16), .ZN(new_n236));
  INV_X1    g035(.A(G22gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G15gat), .ZN(new_n238));
  INV_X1    g037(.A(G15gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G22gat), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT96), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT96), .B1(new_n238), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n236), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT97), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT96), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n239), .A2(G22gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n237), .A2(G15gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT96), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n235), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n245), .A2(new_n252), .A3(G8gat), .ZN(new_n253));
  INV_X1    g052(.A(G8gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n243), .B(new_n251), .C1(new_n244), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n234), .A2(KEYINPUT98), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT98), .B1(new_n234), .B2(new_n256), .ZN(new_n258));
  OAI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(new_n256), .B2(new_n234), .ZN(new_n259));
  NAND2_X1  g058(.A1(G229gat), .A2(G233gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT13), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT98), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n253), .A2(new_n255), .ZN(new_n264));
  INV_X1    g063(.A(new_n233), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n228), .B2(new_n229), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n234), .A2(KEYINPUT98), .A3(new_n256), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n230), .A2(KEYINPUT17), .A3(new_n233), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n271));
  OAI211_X1 g070(.A(new_n264), .B(new_n270), .C1(new_n266), .C2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n269), .A2(KEYINPUT18), .A3(new_n260), .A4(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n260), .C1(new_n257), .C2(new_n258), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT99), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT99), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n269), .A2(new_n277), .A3(new_n260), .A4(new_n272), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G141gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G197gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT11), .B(G169gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT12), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n274), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n274), .B2(new_n280), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(KEYINPUT77), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT77), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n293), .B(new_n294), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n292), .ZN(new_n305));
  OAI221_X1 g104(.A(new_n304), .B1(new_n305), .B2(new_n291), .C1(new_n299), .C2(KEYINPUT78), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT79), .B(G155gat), .Z(new_n307));
  XOR2_X1   g106(.A(KEYINPUT80), .B(G162gat), .Z(new_n308));
  AOI21_X1  g107(.A(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  OAI211_X1 g113(.A(KEYINPUT69), .B(G134gat), .C1(new_n314), .C2(KEYINPUT1), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n316), .B(new_n317), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G127gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n315), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n315), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n315), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G127gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n315), .A2(new_n322), .A3(new_n323), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n290), .B1(new_n312), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n324), .A2(new_n325), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT82), .B1(new_n333), .B2(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n329), .ZN(new_n335));
  INV_X1    g134(.A(new_n310), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT4), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n338), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n336), .B1(new_n326), .B2(new_n330), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n290), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(KEYINPUT5), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n343), .A2(new_n339), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT84), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n351), .A4(new_n339), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n347), .B(new_n332), .C1(new_n348), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n354), .A3(new_n360), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n361), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G8gat), .B(G36gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT74), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  XNOR2_X1  g171(.A(G197gat), .B(G204gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT22), .ZN(new_n374));
  INV_X1    g173(.A(G211gat), .ZN(new_n375));
  INV_X1    g174(.A(G218gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n373), .A3(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(KEYINPUT72), .Z(new_n386));
  INV_X1    g185(.A(G183gat), .ZN(new_n387));
  INV_X1    g186(.A(G190gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT24), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT24), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(KEYINPUT65), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G183gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n396), .B2(G190gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n398), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n399));
  INV_X1    g198(.A(G169gat), .ZN(new_n400));
  INV_X1    g199(.A(G176gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n404), .B2(KEYINPUT23), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n397), .A2(KEYINPUT25), .A3(new_n399), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n399), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n389), .A2(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(new_n409), .B2(KEYINPUT25), .ZN(new_n410));
  AND2_X1   g209(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n411));
  NOR2_X1   g210(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n398), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT68), .B(new_n398), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n398), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n402), .B1(KEYINPUT26), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n387), .B2(new_n388), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  AOI21_X1  g221(.A(G190gat), .B1(new_n422), .B2(G183gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n387), .A2(KEYINPUT27), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n423), .A2(KEYINPUT28), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT27), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT66), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n393), .A2(new_n395), .A3(new_n428), .A4(KEYINPUT27), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT28), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n410), .B1(new_n421), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n386), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n417), .A2(new_n419), .B1(G183gat), .B2(G190gat), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n430), .A2(new_n431), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n425), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n385), .B1(new_n438), .B2(new_n410), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n372), .B(new_n384), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n386), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n438), .B2(new_n410), .ZN(new_n442));
  INV_X1    g241(.A(new_n385), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n383), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n433), .A2(new_n443), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n442), .B2(new_n386), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n372), .B1(new_n447), .B2(new_n384), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n371), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT75), .B(new_n371), .C1(new_n445), .C2(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n434), .ZN(new_n454));
  INV_X1    g253(.A(new_n386), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n454), .A2(new_n455), .B1(new_n443), .B2(new_n433), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT73), .B1(new_n456), .B2(new_n383), .ZN(new_n457));
  INV_X1    g256(.A(new_n371), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n444), .A3(new_n440), .A4(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT30), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n453), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT89), .B1(new_n367), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n464), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n365), .A2(new_n366), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n453), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT31), .B(G50gat), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT29), .B1(new_n381), .B2(new_n382), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n311), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n310), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n303), .B(new_n311), .C1(new_n306), .C2(new_n309), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n383), .B1(new_n480), .B2(new_n434), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n311), .B1(new_n474), .B2(KEYINPUT86), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n310), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n473), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G22gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n492));
  INV_X1    g291(.A(new_n473), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n311), .A3(new_n484), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n481), .B1(new_n495), .B2(new_n310), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n492), .B(new_n493), .C1(new_n496), .C2(new_n479), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n491), .B1(new_n489), .B2(new_n497), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n433), .A2(new_n335), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n438), .A2(new_n410), .A3(new_n333), .ZN(new_n502));
  INV_X1    g301(.A(G227gat), .ZN(new_n503));
  INV_X1    g302(.A(G233gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G43gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n506), .B2(KEYINPUT32), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n506), .B(KEYINPUT32), .C1(new_n507), .C2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT34), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT34), .B(new_n505), .C1(new_n501), .C2(new_n502), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n523), .A3(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT71), .A3(new_n526), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n518), .A2(KEYINPUT71), .A3(new_n524), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n500), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n466), .A2(new_n472), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n498), .A2(new_n499), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n526), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n516), .B2(new_n517), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n532), .A4(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n469), .A2(new_n470), .A3(new_n453), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT35), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n532), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT36), .A3(new_n526), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n453), .A2(new_n462), .A3(new_n464), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT40), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n312), .A2(new_n331), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n348), .B2(new_n353), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n290), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n360), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n343), .A2(new_n290), .A3(new_n344), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT39), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n550), .B2(new_n290), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n548), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n290), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT39), .A3(new_n554), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(KEYINPUT40), .A3(new_n360), .A4(new_n552), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n560), .A3(new_n362), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n532), .B1(new_n547), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n457), .A2(new_n563), .A3(new_n444), .A4(new_n440), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n447), .B2(new_n383), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n384), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT38), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n567), .A3(new_n371), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n365), .A2(new_n568), .A3(new_n366), .A4(new_n459), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT37), .B1(new_n445), .B2(new_n448), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n564), .A3(new_n371), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT38), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n571), .B2(KEYINPUT38), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n542), .B(new_n546), .C1(new_n562), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n288), .B1(new_n540), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  OR2_X1    g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n580), .B(new_n579), .C1(new_n585), .C2(new_n582), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n588));
  AND2_X1   g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n323), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(KEYINPUT101), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n586), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n256), .B1(KEYINPUT21), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT7), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(G85gat), .A3(G92gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n616), .A2(new_n620), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n270), .B(new_n624), .C1(new_n266), .C2(new_n271), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n234), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n610), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n610), .A3(new_n628), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n630), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n608), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n587), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n623), .B(new_n622), .C1(new_n593), .C2(KEYINPUT102), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n623), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n592), .B2(new_n595), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n640), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n640), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n650), .A3(new_n645), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n639), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n367), .A2(KEYINPUT104), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n470), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n577), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT105), .B(G1gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n577), .A2(new_n465), .A3(new_n661), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT106), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(G8gat), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n671), .A2(new_n670), .A3(new_n673), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n527), .A2(new_n528), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n577), .A2(new_n239), .A3(new_n678), .A4(new_n661), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n577), .A2(new_n661), .ZN(new_n680));
  INV_X1    g479(.A(new_n546), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n679), .B1(new_n682), .B2(new_n239), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n541), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT107), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n685), .B(new_n687), .ZN(G1327gat));
  AOI21_X1  g487(.A(new_n638), .B1(new_n540), .B2(new_n576), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n288), .A2(new_n608), .A3(new_n660), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n689), .A2(new_n212), .A3(new_n666), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n540), .A2(new_n576), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n637), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n694), .A3(KEYINPUT44), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n666), .A2(new_n697), .A3(new_n698), .A4(new_n690), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n692), .B1(new_n699), .B2(new_n212), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1328gat));
  AND2_X1   g501(.A1(new_n689), .A2(new_n690), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n213), .A3(new_n465), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n465), .A2(new_n697), .A3(new_n698), .A4(new_n690), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n213), .B2(new_n707), .ZN(G1329gat));
  NAND4_X1  g507(.A1(new_n697), .A2(new_n681), .A3(new_n698), .A4(new_n690), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(new_n206), .A3(new_n678), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT47), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  AOI211_X1 g514(.A(KEYINPUT111), .B(new_n715), .C1(new_n710), .C2(new_n711), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n716), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n703), .A2(new_n203), .A3(new_n541), .ZN(new_n718));
  AND4_X1   g517(.A1(new_n541), .A2(new_n697), .A3(new_n698), .A4(new_n690), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n203), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1331gat));
  INV_X1    g521(.A(new_n288), .ZN(new_n723));
  INV_X1    g522(.A(new_n660), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n723), .A2(new_n639), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n693), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n666), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g528(.A1(new_n726), .A2(KEYINPUT112), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(KEYINPUT112), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n465), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT49), .B(G64gat), .Z(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n681), .A3(new_n731), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G71gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  INV_X1    g538(.A(G71gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n727), .B2(new_n678), .ZN(new_n742));
  INV_X1    g541(.A(new_n678), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n726), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n738), .A2(new_n739), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n739), .B1(new_n738), .B2(new_n745), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n541), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n723), .A2(new_n608), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n724), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n697), .A2(new_n698), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n665), .ZN(new_n755));
  INV_X1    g554(.A(new_n689), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n756), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT51), .B1(new_n756), .B2(new_n752), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n660), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n666), .A2(new_n611), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  OAI21_X1  g560(.A(G92gat), .B1(new_n754), .B2(new_n547), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n465), .A2(new_n612), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n762), .B(new_n766), .C1(new_n759), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1337gat));
  NOR2_X1   g567(.A1(new_n754), .A2(new_n546), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(G99gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n678), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n769), .A2(new_n770), .B1(new_n759), .B2(new_n771), .ZN(G1338gat));
  OAI21_X1  g571(.A(G106gat), .B1(new_n754), .B2(new_n532), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n532), .A2(G106gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n660), .A3(new_n758), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT115), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT115), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1339gat));
  NOR3_X1   g579(.A1(new_n723), .A2(new_n639), .A3(new_n660), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  INV_X1    g581(.A(new_n260), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n272), .B1(new_n257), .B2(new_n258), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n234), .A2(new_n256), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n267), .B2(new_n268), .ZN(new_n786));
  INV_X1    g585(.A(new_n261), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n783), .A2(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n284), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n259), .A2(new_n261), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n260), .B1(new_n269), .B2(new_n272), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT117), .B(new_n284), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n274), .A2(new_n280), .A3(new_n285), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n660), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(new_n640), .C1(new_n646), .C2(new_n648), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n656), .ZN(new_n799));
  INV_X1    g598(.A(new_n648), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n644), .A2(new_n645), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n800), .B(new_n650), .C1(new_n801), .C2(new_n642), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n649), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n657), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n285), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n262), .A2(new_n273), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n815), .B2(new_n795), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n638), .B1(new_n796), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n637), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n794), .A2(new_n795), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n608), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n781), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n541), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n547), .A3(new_n678), .A4(new_n666), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n318), .A3(new_n288), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n825), .A2(new_n465), .A3(new_n537), .A4(new_n665), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n723), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n828), .A2(new_n830), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n827), .B2(new_n724), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n660), .A2(new_n320), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT118), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1341gat));
  XOR2_X1   g635(.A(KEYINPUT69), .B(G127gat), .Z(new_n837));
  NOR3_X1   g636(.A1(new_n827), .A2(new_n824), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n829), .A2(new_n608), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT119), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n840), .B2(new_n837), .ZN(G1342gat));
  NAND3_X1  g640(.A1(new_n829), .A2(new_n317), .A3(new_n637), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n827), .B2(new_n638), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n681), .A2(new_n665), .A3(new_n465), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n532), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n817), .A2(KEYINPUT120), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n818), .B1(new_n286), .B2(new_n287), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n794), .A2(new_n795), .A3(new_n660), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n637), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n822), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n824), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n661), .A2(new_n288), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n850), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n824), .B1(new_n854), .B2(new_n821), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n532), .B1(new_n860), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n847), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n288), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n546), .A2(new_n541), .ZN(new_n865));
  NOR4_X1   g664(.A1(new_n825), .A2(new_n465), .A3(new_n665), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n295), .A3(new_n723), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(G148gat), .C1(new_n863), .C2(new_n724), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT121), .B(new_n848), .C1(new_n825), .C2(new_n532), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n858), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n849), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n847), .A2(new_n660), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G148gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n872), .B1(new_n881), .B2(KEYINPUT59), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n297), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(KEYINPUT122), .A3(new_n870), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n871), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n297), .A3(new_n660), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1345gat));
  OAI21_X1  g686(.A(new_n307), .B1(new_n863), .B2(new_n824), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n824), .A2(new_n307), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1346gat));
  NOR2_X1   g690(.A1(new_n638), .A2(new_n308), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n866), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT123), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n308), .B1(new_n863), .B2(new_n638), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n665), .A2(new_n465), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT126), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT126), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n826), .A2(new_n678), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n400), .A3(new_n288), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n825), .A2(new_n666), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT124), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n537), .A2(new_n547), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT125), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n723), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n901), .B1(new_n906), .B2(new_n400), .ZN(G1348gat));
  OAI21_X1  g706(.A(G176gat), .B1(new_n900), .B2(new_n724), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n903), .A2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n660), .A2(new_n401), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(G1349gat));
  OAI21_X1  g712(.A(new_n396), .B1(new_n900), .B2(new_n824), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n422), .A2(G183gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n608), .A2(new_n915), .A3(new_n424), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g717(.A1(new_n900), .A2(new_n638), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(G190gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(G190gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n637), .A2(new_n388), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n921), .A2(new_n922), .B1(new_n909), .B2(new_n923), .ZN(G1351gat));
  NOR2_X1   g723(.A1(new_n865), .A2(new_n547), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n903), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n723), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n898), .A2(new_n546), .A3(new_n899), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n878), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n723), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n660), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n926), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT62), .B1(new_n926), .B2(new_n934), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n930), .A2(new_n660), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n935), .B(new_n936), .C1(new_n933), .C2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n375), .A3(new_n608), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n608), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n376), .A3(new_n637), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n930), .A2(new_n637), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n376), .ZN(G1355gat));
endmodule


