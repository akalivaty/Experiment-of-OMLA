//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n191), .A2(new_n193), .B1(G143), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT66), .B(new_n189), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(G146), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n194), .A2(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n188), .A2(G128), .A3(new_n191), .A4(new_n193), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n197), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n209), .B2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n210), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n208), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n210), .A3(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n194), .A2(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n198), .A2(G146), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT0), .A4(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n188), .A2(new_n230), .A3(KEYINPUT0), .A4(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n188), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n237), .A2(KEYINPUT67), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n249), .A3(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n222), .A2(new_n236), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n234), .B1(new_n229), .B2(new_n231), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n225), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n222), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n250), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT30), .B1(new_n222), .B2(new_n236), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT29), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n253), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT68), .B1(new_n241), .B2(new_n249), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n236), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n226), .A2(new_n227), .A3(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n191), .A2(new_n193), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n201), .A2(new_n205), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(KEYINPUT66), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n220), .B1(new_n277), .B2(new_n206), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n250), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n222), .B2(new_n236), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT28), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n272), .B2(new_n278), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT71), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n255), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n282), .A2(new_n285), .A3(new_n267), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT29), .A4(new_n267), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT72), .B1(new_n272), .B2(new_n278), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n252), .A2(new_n253), .B1(new_n257), .B2(new_n225), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n222), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n270), .A2(new_n271), .ZN(new_n297));
  INV_X1    g111(.A(new_n236), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n278), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT28), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n292), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G472), .B1(new_n291), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n208), .A2(new_n221), .B1(new_n225), .B2(new_n257), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n259), .B(new_n250), .C1(KEYINPUT30), .C2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n255), .A3(new_n267), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n256), .B1(new_n278), .B2(new_n298), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n280), .B1(new_n222), .B2(new_n258), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n279), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(KEYINPUT70), .A3(new_n267), .A4(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n282), .A2(new_n285), .A3(new_n287), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n308), .A2(new_n255), .A3(new_n267), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n268), .B1(KEYINPUT31), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(G472), .A2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT32), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n187), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G472), .ZN(new_n330));
  INV_X1    g144(.A(new_n292), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n300), .A2(KEYINPUT73), .A3(KEYINPUT28), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT73), .B1(new_n300), .B2(KEYINPUT28), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n269), .B2(new_n288), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n325), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n317), .B2(new_n320), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n312), .A2(new_n316), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n319), .A2(KEYINPUT31), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n250), .B1(new_n278), .B2(new_n298), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n283), .B1(new_n342), .B2(new_n255), .ZN(new_n343));
  AOI211_X1 g157(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n294), .C2(new_n222), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n286), .B1(new_n255), .B2(new_n283), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n341), .B1(new_n346), .B2(new_n267), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n322), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n324), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n339), .A2(new_n349), .A3(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n329), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n290), .ZN(new_n353));
  OR2_X1    g167(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT23), .B1(new_n196), .B2(G119), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n196), .A2(G119), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT75), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT75), .B1(new_n242), .B2(G128), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n242), .A2(G128), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT23), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT76), .B1(new_n361), .B2(G110), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n356), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT24), .B(G110), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n366));
  INV_X1    g180(.A(G110), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n357), .A2(new_n360), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G125), .ZN(new_n371));
  INV_X1    g185(.A(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT16), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n370), .A3(G125), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  MUX2_X1   g191(.A(new_n374), .B(new_n377), .S(G146), .Z(new_n378));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n377), .A2(new_n194), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n194), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n363), .A2(new_n364), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n361), .B2(G110), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G137), .ZN(new_n386));
  INV_X1    g200(.A(G953), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G221), .A3(G234), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n379), .B2(new_n385), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n354), .B1(new_n393), .B2(new_n290), .ZN(new_n394));
  NOR2_X1   g208(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n395));
  NOR4_X1   g209(.A1(new_n391), .A2(new_n392), .A3(G902), .A4(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n353), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n353), .A2(G902), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT78), .Z(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n208), .A2(new_n372), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n257), .A2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G224), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n242), .A3(G116), .ZN(new_n411));
  OAI211_X1 g225(.A(G113), .B(new_n411), .C1(new_n246), .C2(new_n410), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n247), .B2(new_n246), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT79), .B(G101), .ZN(new_n414));
  INV_X1    g228(.A(G104), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT3), .B1(new_n415), .B2(G107), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n417));
  INV_X1    g231(.A(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G104), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(G107), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n414), .A2(new_n416), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(G104), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n420), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G101), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n413), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G101), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n421), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT80), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n431), .A3(new_n421), .A4(KEYINPUT4), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n427), .A2(new_n434), .A3(G101), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n250), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n426), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT83), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n430), .B2(new_n432), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  NOR4_X1   g257(.A1(new_n441), .A2(new_n442), .A3(new_n426), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n437), .ZN(new_n445));
  INV_X1    g259(.A(new_n426), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n440), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n446), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT6), .A4(new_n443), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n450), .B(new_n443), .C1(new_n441), .C2(new_n426), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n409), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n442), .B1(new_n449), .B2(new_n443), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n439), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n407), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n405), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n439), .B(KEYINPUT8), .Z(new_n463));
  NAND2_X1  g277(.A1(new_n413), .A2(new_n425), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n446), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n460), .B1(new_n407), .B2(KEYINPUT85), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT85), .B2(new_n407), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n403), .B2(new_n404), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n462), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n459), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n456), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n456), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n402), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(G475), .A2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n371), .A2(new_n373), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n194), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n374), .B2(G146), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n374), .A2(new_n481), .A3(G146), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT18), .A2(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n263), .A2(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n198), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT18), .A3(G131), .A4(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT88), .B1(new_n477), .B2(new_n194), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n479), .A3(new_n478), .A4(new_n483), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n492), .A2(new_n218), .A3(new_n487), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n374), .B(KEYINPUT19), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n380), .B(new_n500), .C1(G146), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n415), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n508), .A3(new_n499), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT17), .B(G131), .C1(new_n488), .C2(new_n489), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n509), .A2(new_n380), .A3(new_n381), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n497), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n476), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n514));
  OAI21_X1  g328(.A(KEYINPUT89), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n497), .A2(new_n511), .A3(new_n505), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n505), .B1(new_n497), .B2(new_n502), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n475), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  INV_X1    g333(.A(new_n514), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(new_n475), .C1(new_n516), .C2(new_n517), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n507), .A2(new_n512), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT90), .A3(new_n522), .A4(new_n475), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n515), .A2(new_n521), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n505), .B1(new_n497), .B2(new_n511), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n290), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT91), .B(new_n290), .C1(new_n516), .C2(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(G475), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT9), .B(G234), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n352), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G128), .B(G143), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n209), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n244), .B2(G122), .ZN(new_n542));
  INV_X1    g356(.A(G122), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT92), .A3(G116), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n244), .A2(G122), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n418), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n546), .B(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n418), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n546), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G107), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT13), .B1(new_n196), .B2(G143), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n209), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n556), .A2(new_n539), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n539), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n554), .A2(new_n547), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n538), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n550), .A2(new_n545), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n547), .B(new_n540), .C1(new_n561), .C2(new_n418), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n554), .A2(new_n547), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n558), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n565), .A3(new_n537), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n566), .A3(KEYINPUT93), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(new_n538), .C1(new_n552), .C2(new_n559), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n290), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(new_n290), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n387), .A2(G952), .ZN(new_n577));
  INV_X1    g391(.A(G234), .ZN(new_n578));
  INV_X1    g392(.A(G237), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n290), .B(new_n387), .C1(G234), .C2(G237), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n535), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G469), .ZN(new_n587));
  INV_X1    g401(.A(new_n225), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n197), .A2(new_n425), .A3(new_n206), .A4(new_n207), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n188), .B2(G128), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n421), .B(new_n424), .C1(new_n275), .C2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n588), .B2(KEYINPUT82), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n593), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n592), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n433), .A2(new_n257), .A3(new_n435), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n425), .A2(new_n597), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n208), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n588), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(G110), .B(G140), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n387), .A2(G227), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n596), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n592), .A2(new_n600), .A3(new_n597), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n600), .B1(new_n592), .B2(new_n597), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n605), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n257), .A2(new_n435), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n432), .B2(new_n430), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n225), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n610), .B1(new_n617), .B2(new_n606), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n587), .B(new_n290), .C1(new_n611), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(G469), .A2(G902), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n596), .A2(new_n606), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n609), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n606), .A3(new_n610), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(G469), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G221), .B1(new_n536), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n474), .A2(new_n586), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n351), .A2(new_n401), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT94), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n414), .ZN(G3));
  AND2_X1   g445(.A1(new_n570), .A2(new_n571), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n560), .A2(KEYINPUT33), .A3(new_n566), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n567), .A2(new_n634), .A3(new_n569), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n567), .A2(KEYINPUT97), .A3(new_n634), .A4(new_n569), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n571), .A2(G902), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n632), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n535), .A2(new_n641), .A3(new_n584), .ZN(new_n642));
  INV_X1    g456(.A(new_n471), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n452), .B(KEYINPUT6), .ZN(new_n644));
  INV_X1    g458(.A(new_n447), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n457), .A2(new_n645), .A3(new_n458), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n408), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n469), .B1(new_n440), .B2(new_n444), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n290), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n643), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n456), .A2(new_n470), .A3(new_n471), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n402), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n473), .B2(KEYINPUT96), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n642), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n401), .A2(new_n625), .A3(new_n626), .ZN(new_n657));
  NAND2_X1  g471(.A1(KEYINPUT95), .A2(G472), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AOI211_X1 g473(.A(G902), .B(new_n659), .C1(new_n317), .C2(new_n320), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n321), .B2(new_n290), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n655), .A2(new_n653), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n515), .B(new_n521), .C1(new_n520), .C2(new_n518), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n534), .A3(new_n576), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(new_n584), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n662), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n472), .A2(new_n473), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n627), .A3(new_n654), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n379), .A2(new_n385), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT36), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n389), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n676), .B(new_n678), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n399), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n397), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n534), .A3(new_n528), .A4(new_n585), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n661), .A3(new_n660), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  AOI21_X1  g500(.A(new_n666), .B1(new_n329), .B2(new_n350), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n625), .A2(new_n626), .A3(new_n681), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n582), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n580), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n688), .A2(new_n668), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT98), .B(G128), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G30));
  XOR2_X1   g510(.A(new_n691), .B(KEYINPUT39), .Z(new_n697));
  OR2_X1    g511(.A1(new_n627), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n300), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n319), .B1(new_n701), .B2(new_n267), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n330), .B1(new_n702), .B2(new_n290), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n338), .A2(new_n703), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n704), .A2(KEYINPUT99), .A3(new_n328), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT99), .B1(new_n704), .B2(new_n328), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n674), .B(KEYINPUT38), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n528), .A2(new_n534), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n576), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n710), .A2(new_n654), .A3(new_n681), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n707), .A3(new_n708), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  AND2_X1   g527(.A1(new_n655), .A2(new_n653), .ZN(new_n714));
  INV_X1    g528(.A(new_n640), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n633), .B(new_n715), .C1(new_n637), .C2(new_n638), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n709), .B(new_n691), .C1(new_n632), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n688), .A2(new_n717), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n328), .A2(new_n336), .A3(new_n338), .A4(new_n187), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT74), .B1(new_n339), .B2(new_n349), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n714), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n351), .A2(KEYINPUT100), .A3(new_n714), .A4(new_n718), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n619), .A2(new_n727), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n599), .A2(new_n601), .B1(new_n208), .B2(new_n604), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n588), .B1(new_n729), .B2(new_n603), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n614), .A2(new_n225), .A3(new_n616), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n609), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n596), .A2(new_n606), .A3(new_n610), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n587), .B1(new_n734), .B2(new_n290), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n727), .B(new_n587), .C1(new_n734), .C2(new_n290), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n626), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n351), .A2(new_n656), .A3(new_n401), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n351), .A2(new_n401), .A3(new_n670), .A4(new_n739), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NOR2_X1   g558(.A1(new_n738), .A2(new_n682), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n687), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  AOI21_X1  g561(.A(new_n330), .B1(new_n321), .B2(new_n290), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n345), .A2(new_n344), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n332), .B2(new_n333), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(new_n268), .B1(KEYINPUT31), .B2(new_n319), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n340), .B1(new_n751), .B2(KEYINPUT103), .ZN(new_n752));
  INV_X1    g566(.A(new_n749), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n303), .B2(new_n304), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n341), .B1(new_n754), .B2(new_n267), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n322), .B(KEYINPUT102), .Z(new_n759));
  AOI21_X1  g573(.A(new_n748), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n738), .A2(new_n666), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n710), .A2(new_n584), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n401), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  INV_X1    g578(.A(new_n759), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n752), .B2(new_n757), .ZN(new_n766));
  INV_X1    g580(.A(new_n681), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n766), .A2(new_n767), .A3(new_n748), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n738), .A2(new_n666), .A3(new_n717), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  NAND2_X1  g585(.A1(new_n328), .A2(KEYINPUT105), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n323), .B1(new_n317), .B2(new_n320), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(KEYINPUT32), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n326), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n772), .A2(KEYINPUT106), .A3(new_n326), .A4(new_n775), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n306), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n717), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n472), .A2(new_n473), .A3(new_n654), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n619), .A2(KEYINPUT104), .A3(new_n624), .A4(new_n620), .ZN(new_n783));
  INV_X1    g597(.A(new_n626), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT104), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n625), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n780), .A2(new_n789), .A3(new_n401), .ZN(new_n790));
  INV_X1    g604(.A(new_n401), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n329), .B2(new_n350), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n782), .A2(new_n786), .A3(new_n783), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n781), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n790), .B1(new_n794), .B2(KEYINPUT42), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NOR2_X1   g610(.A1(new_n668), .A2(new_n692), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n351), .A2(new_n401), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT107), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n792), .A2(new_n800), .A3(new_n797), .A4(new_n793), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND2_X1  g617(.A1(new_n622), .A2(new_n623), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n587), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n622), .A2(KEYINPUT45), .A3(new_n623), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n620), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT46), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT46), .A3(new_n620), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n619), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n626), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n697), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n641), .A2(new_n709), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT43), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT110), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(KEYINPUT110), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n820), .A2(KEYINPUT43), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT109), .B1(new_n820), .B2(KEYINPUT43), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n822), .A2(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n681), .B1(new_n661), .B2(new_n660), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n819), .B1(new_n830), .B2(KEYINPUT44), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n650), .A2(new_n652), .A3(new_n402), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n830), .B2(KEYINPUT44), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT44), .ZN(new_n834));
  OAI211_X1 g648(.A(KEYINPUT111), .B(new_n834), .C1(new_n828), .C2(new_n829), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n818), .A2(new_n831), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n216), .ZN(G39));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT47), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n626), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT112), .B1(new_n816), .B2(new_n626), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n839), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n626), .ZN(new_n846));
  NAND2_X1  g660(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n351), .A2(new_n401), .A3(new_n717), .A4(new_n832), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  INV_X1    g666(.A(new_n736), .ZN(new_n853));
  INV_X1    g667(.A(new_n737), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT49), .Z(new_n856));
  NAND4_X1  g670(.A1(new_n820), .A2(new_n401), .A3(new_n626), .A4(new_n402), .ZN(new_n857));
  OR4_X1    g671(.A1(new_n707), .A2(new_n856), .A3(new_n708), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  INV_X1    g673(.A(new_n707), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n738), .A2(new_n832), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n791), .A2(new_n580), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n709), .A2(new_n716), .A3(new_n632), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n822), .A2(new_n823), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n826), .A2(new_n827), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n580), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n317), .B1(new_n755), .B2(new_n756), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n759), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n748), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n681), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n864), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n708), .A2(new_n402), .A3(new_n738), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n766), .A2(new_n791), .A3(new_n748), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n867), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n867), .A2(new_n875), .A3(KEYINPUT50), .A4(new_n876), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n859), .B1(new_n881), .B2(KEYINPUT120), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n784), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n842), .A2(new_n848), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n867), .A2(new_n876), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n832), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n879), .A2(new_n880), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n867), .A2(new_n861), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n768), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n892), .A3(new_n864), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n882), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n780), .A2(new_n401), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT48), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n709), .B1(new_n632), .B2(new_n716), .ZN(new_n901));
  INV_X1    g715(.A(new_n761), .ZN(new_n902));
  OAI221_X1 g716(.A(new_n577), .B1(new_n900), .B2(new_n901), .C1(new_n887), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n893), .B1(new_n886), .B2(new_n888), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n896), .B(new_n904), .C1(KEYINPUT51), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n768), .A2(new_n769), .B1(new_n687), .B2(new_n693), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n681), .A2(new_n692), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT115), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n786), .A2(new_n783), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n666), .A2(new_n710), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n707), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n725), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n725), .A2(new_n916), .A3(new_n908), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n763), .A2(new_n740), .A3(new_n743), .ZN(new_n919));
  INV_X1    g733(.A(new_n584), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n402), .C1(new_n472), .C2(new_n473), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n528), .A2(new_n534), .A3(new_n576), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT114), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n901), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n709), .B(new_n923), .C1(new_n632), .C2(new_n716), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n927), .A2(new_n662), .B1(new_n675), .B2(new_n683), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n746), .A2(new_n928), .A3(new_n629), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n919), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n576), .A2(new_n692), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n667), .A3(new_n534), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n688), .A2(new_n832), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n720), .B2(new_n719), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n873), .B2(new_n787), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n799), .B2(new_n801), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n795), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n907), .B1(new_n918), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n930), .A2(new_n795), .A3(new_n936), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n914), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(KEYINPUT53), .A3(new_n917), .A4(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(KEYINPUT118), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n917), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT117), .B(new_n907), .C1(new_n946), .C2(new_n937), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n939), .A2(KEYINPUT53), .A3(new_n917), .A4(new_n915), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n936), .A2(new_n795), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(new_n930), .A3(new_n941), .A4(new_n917), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT117), .B1(new_n951), .B2(new_n907), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT54), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n955), .B(KEYINPUT54), .C1(new_n949), .C2(new_n952), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n906), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n858), .B1(new_n957), .B2(new_n958), .ZN(G75));
  NOR2_X1   g773(.A1(new_n387), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n290), .B1(new_n938), .B2(new_n942), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT56), .B1(new_n962), .B2(G210), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n448), .A2(new_n455), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n408), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n456), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT55), .Z(new_n967));
  OAI21_X1  g781(.A(new_n961), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n967), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n963), .A2(KEYINPUT121), .A3(new_n967), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G51));
  NAND2_X1  g787(.A1(new_n938), .A2(new_n942), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n943), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n620), .B(KEYINPUT57), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n734), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(G902), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(new_n811), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n960), .B1(new_n977), .B2(new_n979), .ZN(G54));
  AND3_X1   g794(.A1(new_n962), .A2(KEYINPUT58), .A3(G475), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n961), .B1(new_n981), .B2(new_n526), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n526), .B2(new_n981), .ZN(G60));
  NAND2_X1  g797(.A1(G478), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT59), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n639), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n961), .B1(new_n975), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n639), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n954), .A2(new_n956), .A3(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(G63));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT122), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n974), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n393), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n974), .A2(new_n679), .A3(new_n994), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n961), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G66));
  OAI21_X1  g815(.A(G953), .B1(new_n583), .B2(new_n406), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n930), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n964), .B1(G898), .B2(new_n387), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  AOI21_X1  g819(.A(new_n387), .B1(G227), .B2(G900), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n313), .A2(new_n259), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n501), .B(KEYINPUT123), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(G900), .B2(G953), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n836), .B1(new_n849), .B2(new_n850), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n818), .A2(new_n897), .A3(new_n912), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n725), .A2(new_n908), .ZN(new_n1013));
  AND4_X1   g827(.A1(new_n795), .A2(new_n1012), .A3(new_n802), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1010), .B1(new_n1015), .B2(G953), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1009), .B(KEYINPUT124), .Z(new_n1018));
  NAND3_X1  g832(.A1(new_n712), .A2(new_n725), .A3(new_n908), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT125), .Z(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n832), .B(new_n698), .C1(new_n925), .C2(new_n926), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n792), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1021), .A2(new_n1011), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1018), .B1(new_n1025), .B2(new_n387), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1006), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1006), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1025), .A2(new_n387), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1028), .B(new_n1016), .C1(new_n1029), .C2(new_n1018), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  INV_X1    g847(.A(new_n930), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1033), .B1(new_n1015), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n315), .B(KEYINPUT126), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n268), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT127), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n960), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1033), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1036), .A2(new_n268), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n319), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n315), .A2(new_n267), .ZN(new_n1044));
  OAI221_X1 g858(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .C1(new_n949), .C2(new_n952), .ZN(new_n1045));
  AND3_X1   g859(.A1(new_n1039), .A2(new_n1042), .A3(new_n1045), .ZN(G57));
endmodule


