

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758;

  INV_X1 U373 ( .A(n726), .ZN(n353) );
  NOR2_X1 U374 ( .A1(n664), .A2(n359), .ZN(n393) );
  NOR2_X1 U375 ( .A1(n532), .A2(n560), .ZN(n654) );
  XNOR2_X1 U376 ( .A(n386), .B(G134), .ZN(n529) );
  XNOR2_X1 U377 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n492) );
  INV_X1 U378 ( .A(n352), .ZN(n716) );
  NAND2_X1 U379 ( .A1(n354), .A2(n353), .ZN(n352) );
  XNOR2_X1 U380 ( .A(n714), .B(n355), .ZN(n354) );
  INV_X1 U381 ( .A(n713), .ZN(n355) );
  XNOR2_X2 U382 ( .A(n567), .B(n566), .ZN(n633) );
  XNOR2_X2 U383 ( .A(n743), .B(n477), .ZN(n615) );
  XNOR2_X1 U384 ( .A(G146), .B(KEYINPUT67), .ZN(n416) );
  AND2_X1 U385 ( .A1(n404), .A2(n403), .ZN(n611) );
  NAND2_X1 U386 ( .A1(n532), .A2(n560), .ZN(n660) );
  NOR2_X2 U387 ( .A1(n607), .A2(n587), .ZN(n589) );
  NOR2_X1 U388 ( .A1(n607), .A2(n703), .ZN(n585) );
  AND2_X2 U389 ( .A1(n389), .A2(n391), .ZN(n369) );
  XNOR2_X2 U390 ( .A(n486), .B(n485), .ZN(n549) );
  NOR2_X2 U391 ( .A1(n756), .A2(n633), .ZN(n568) );
  XNOR2_X2 U392 ( .A(n434), .B(KEYINPUT35), .ZN(n755) );
  XNOR2_X2 U393 ( .A(n501), .B(n500), .ZN(n557) );
  NAND2_X1 U394 ( .A1(n600), .A2(n678), .ZN(n687) );
  XNOR2_X1 U395 ( .A(n416), .B(G131), .ZN(n518) );
  BUF_X1 U396 ( .A(n734), .Z(n356) );
  XNOR2_X2 U397 ( .A(n395), .B(KEYINPUT39), .ZN(n575) );
  NOR2_X1 U398 ( .A1(n548), .A2(n600), .ZN(n464) );
  INV_X1 U399 ( .A(G237), .ZN(n499) );
  XNOR2_X1 U400 ( .A(n467), .B(n518), .ZN(n415) );
  XNOR2_X1 U401 ( .A(KEYINPUT68), .B(G137), .ZN(n466) );
  INV_X1 U402 ( .A(G902), .ZN(n457) );
  AND2_X1 U403 ( .A1(n674), .A2(n429), .ZN(n428) );
  XNOR2_X1 U404 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U405 ( .A(KEYINPUT5), .B(G119), .ZN(n471) );
  XNOR2_X1 U406 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n470) );
  XNOR2_X1 U407 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n469) );
  INV_X1 U408 ( .A(n757), .ZN(n412) );
  XNOR2_X1 U409 ( .A(n433), .B(n432), .ZN(n488) );
  XNOR2_X1 U410 ( .A(G116), .B(G113), .ZN(n432) );
  XNOR2_X1 U411 ( .A(n468), .B(G101), .ZN(n433) );
  INV_X1 U412 ( .A(KEYINPUT3), .ZN(n468) );
  NOR2_X1 U413 ( .A1(n401), .A2(n400), .ZN(n403) );
  AND2_X1 U414 ( .A1(n402), .A2(KEYINPUT44), .ZN(n401) );
  NAND2_X1 U415 ( .A1(n362), .A2(n643), .ZN(n400) );
  XNOR2_X1 U416 ( .A(n371), .B(n370), .ZN(n524) );
  INV_X1 U417 ( .A(KEYINPUT8), .ZN(n370) );
  XNOR2_X1 U418 ( .A(G113), .B(G122), .ZN(n512) );
  XNOR2_X1 U419 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U420 ( .A(G107), .B(G104), .Z(n487) );
  XNOR2_X1 U421 ( .A(n494), .B(n493), .ZN(n495) );
  INV_X1 U422 ( .A(n492), .ZN(n493) );
  INV_X1 U423 ( .A(G128), .ZN(n465) );
  NAND2_X1 U424 ( .A1(n378), .A2(n377), .ZN(n376) );
  AND2_X1 U425 ( .A1(n591), .A2(KEYINPUT28), .ZN(n377) );
  AND2_X1 U426 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U427 ( .A(n407), .B(n491), .ZN(n735) );
  XNOR2_X1 U428 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U429 ( .A(n488), .B(n487), .ZN(n407) );
  XNOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n489) );
  XOR2_X1 U431 ( .A(G107), .B(KEYINPUT7), .Z(n526) );
  XNOR2_X1 U432 ( .A(G116), .B(G122), .ZN(n528) );
  INV_X1 U433 ( .A(KEYINPUT9), .ZN(n373) );
  NOR2_X1 U434 ( .A1(n657), .A2(n374), .ZN(n542) );
  NAND2_X1 U435 ( .A1(n375), .A2(n378), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n531), .B(G478), .ZN(n560) );
  OR2_X2 U437 ( .A1(n431), .A2(n581), .ZN(n582) );
  OR2_X1 U438 ( .A1(n428), .A2(KEYINPUT47), .ZN(n426) );
  AND2_X1 U439 ( .A1(n425), .A2(n535), .ZN(n424) );
  AND2_X1 U440 ( .A1(n428), .A2(KEYINPUT47), .ZN(n425) );
  OR2_X1 U441 ( .A1(n654), .A2(n533), .ZN(n674) );
  XOR2_X1 U442 ( .A(G122), .B(KEYINPUT16), .Z(n490) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n442) );
  INV_X1 U444 ( .A(n631), .ZN(n363) );
  INV_X1 U445 ( .A(KEYINPUT84), .ZN(n365) );
  XNOR2_X1 U446 ( .A(G128), .B(KEYINPUT24), .ZN(n449) );
  INV_X1 U447 ( .A(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U448 ( .A(KEYINPUT15), .B(G902), .ZN(n612) );
  XNOR2_X1 U449 ( .A(KEYINPUT10), .B(G125), .ZN(n385) );
  XNOR2_X1 U450 ( .A(G143), .B(G104), .ZN(n514) );
  XOR2_X1 U451 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n510) );
  XNOR2_X1 U452 ( .A(G101), .B(G110), .ZN(n483) );
  XNOR2_X1 U453 ( .A(n408), .B(n735), .ZN(n636) );
  XNOR2_X1 U454 ( .A(n410), .B(n409), .ZN(n408) );
  XNOR2_X1 U455 ( .A(n497), .B(n495), .ZN(n410) );
  XNOR2_X1 U456 ( .A(n562), .B(n561), .ZN(n702) );
  XNOR2_X1 U457 ( .A(n589), .B(n588), .ZN(n592) );
  INV_X1 U458 ( .A(KEYINPUT22), .ZN(n588) );
  XNOR2_X1 U459 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U460 ( .A(KEYINPUT103), .ZN(n418) );
  BUF_X1 U461 ( .A(n541), .Z(n683) );
  XNOR2_X1 U462 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U463 ( .A1(n458), .A2(n457), .ZN(n463) );
  XNOR2_X1 U464 ( .A(n527), .B(n372), .ZN(n530) );
  XNOR2_X1 U465 ( .A(n528), .B(n373), .ZN(n372) );
  AND2_X1 U466 ( .A1(n618), .A2(G953), .ZN(n726) );
  XNOR2_X1 U467 ( .A(n574), .B(KEYINPUT102), .ZN(n757) );
  OR2_X1 U468 ( .A1(n571), .A2(n590), .ZN(n572) );
  XNOR2_X1 U469 ( .A(n564), .B(KEYINPUT42), .ZN(n756) );
  NOR2_X1 U470 ( .A1(n702), .A2(n563), .ZN(n564) );
  XNOR2_X1 U471 ( .A(n543), .B(KEYINPUT106), .ZN(n544) );
  NOR2_X1 U472 ( .A1(n539), .A2(n571), .ZN(n545) );
  INV_X1 U473 ( .A(n586), .ZN(n435) );
  AND2_X1 U474 ( .A1(n758), .A2(n406), .ZN(n357) );
  AND2_X1 U475 ( .A1(n393), .A2(n570), .ZN(n358) );
  OR2_X1 U476 ( .A1(n556), .A2(n555), .ZN(n359) );
  XOR2_X1 U477 ( .A(KEYINPUT72), .B(G472), .Z(n360) );
  XOR2_X1 U478 ( .A(n512), .B(n511), .Z(n361) );
  XOR2_X1 U479 ( .A(n609), .B(KEYINPUT99), .Z(n362) );
  NAND2_X1 U480 ( .A1(n464), .A2(n678), .ZN(n540) );
  INV_X1 U481 ( .A(n655), .ZN(n650) );
  INV_X1 U482 ( .A(G140), .ZN(n479) );
  INV_X1 U483 ( .A(KEYINPUT47), .ZN(n430) );
  INV_X1 U484 ( .A(KEYINPUT71), .ZN(n405) );
  AND2_X2 U485 ( .A1(n364), .A2(n363), .ZN(n745) );
  XNOR2_X1 U486 ( .A(n411), .B(n365), .ZN(n364) );
  XNOR2_X1 U487 ( .A(n568), .B(KEYINPUT46), .ZN(n394) );
  NOR2_X1 U488 ( .A1(n537), .A2(n366), .ZN(n538) );
  NAND2_X1 U489 ( .A1(n421), .A2(n423), .ZN(n366) );
  NAND2_X1 U490 ( .A1(n746), .A2(G234), .ZN(n371) );
  XNOR2_X2 U491 ( .A(n367), .B(n360), .ZN(n541) );
  NOR2_X2 U492 ( .A1(n615), .A2(G902), .ZN(n367) );
  NAND2_X1 U493 ( .A1(n745), .A2(n727), .ZN(n666) );
  NAND2_X1 U494 ( .A1(n388), .A2(n358), .ZN(n387) );
  XNOR2_X1 U495 ( .A(n368), .B(n513), .ZN(n520) );
  XNOR2_X1 U496 ( .A(n516), .B(n361), .ZN(n368) );
  NAND2_X1 U497 ( .A1(n655), .A2(n424), .ZN(n423) );
  NOR2_X2 U498 ( .A1(n687), .A2(n686), .ZN(n602) );
  AND2_X1 U499 ( .A1(n597), .A2(KEYINPUT71), .ZN(n397) );
  NAND2_X1 U500 ( .A1(n369), .A2(n387), .ZN(n413) );
  NAND2_X1 U501 ( .A1(n569), .A2(n393), .ZN(n390) );
  INV_X1 U502 ( .A(n598), .ZN(n375) );
  NAND2_X1 U503 ( .A1(n379), .A2(n376), .ZN(n420) );
  INV_X1 U504 ( .A(n540), .ZN(n378) );
  NAND2_X1 U505 ( .A1(n381), .A2(n478), .ZN(n380) );
  INV_X1 U506 ( .A(n591), .ZN(n381) );
  NAND2_X1 U507 ( .A1(n540), .A2(n478), .ZN(n382) );
  NAND2_X1 U508 ( .A1(n383), .A2(n547), .ZN(n556) );
  NAND2_X1 U509 ( .A1(n655), .A2(n384), .ZN(n383) );
  NOR2_X1 U510 ( .A1(n674), .A2(n429), .ZN(n384) );
  NOR2_X4 U511 ( .A1(n563), .A2(n431), .ZN(n655) );
  XNOR2_X2 U512 ( .A(n385), .B(n479), .ZN(n744) );
  XNOR2_X1 U513 ( .A(n386), .B(n498), .ZN(n409) );
  XNOR2_X2 U514 ( .A(n417), .B(n465), .ZN(n386) );
  NAND2_X1 U515 ( .A1(n591), .A2(n670), .ZN(n551) );
  XNOR2_X2 U516 ( .A(n541), .B(KEYINPUT100), .ZN(n591) );
  AND2_X1 U517 ( .A1(n394), .A2(n569), .ZN(n388) );
  NAND2_X1 U518 ( .A1(n390), .A2(n414), .ZN(n389) );
  NAND2_X1 U519 ( .A1(n392), .A2(n414), .ZN(n391) );
  INV_X1 U520 ( .A(n394), .ZN(n392) );
  NAND2_X1 U521 ( .A1(n575), .A2(n654), .ZN(n567) );
  NAND2_X1 U522 ( .A1(n565), .A2(n669), .ZN(n395) );
  NOR2_X2 U523 ( .A1(n552), .A2(n553), .ZN(n565) );
  NAND2_X1 U524 ( .A1(n398), .A2(n396), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n357), .A2(n397), .ZN(n396) );
  NAND2_X1 U526 ( .A1(n399), .A2(n405), .ZN(n398) );
  NAND2_X1 U527 ( .A1(n357), .A2(n597), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n597), .A2(n758), .ZN(n402) );
  INV_X1 U529 ( .A(KEYINPUT44), .ZN(n406) );
  XNOR2_X2 U530 ( .A(n454), .B(G146), .ZN(n497) );
  XNOR2_X1 U531 ( .A(n585), .B(KEYINPUT34), .ZN(n436) );
  XNOR2_X1 U532 ( .A(n448), .B(n447), .ZN(n453) );
  XNOR2_X2 U533 ( .A(n558), .B(KEYINPUT105), .ZN(n673) );
  NAND2_X1 U534 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U535 ( .A(n570), .ZN(n414) );
  XNOR2_X2 U536 ( .A(n529), .B(n415), .ZN(n743) );
  XNOR2_X2 U537 ( .A(KEYINPUT64), .B(G143), .ZN(n417) );
  XNOR2_X2 U538 ( .A(n419), .B(n418), .ZN(n563) );
  NAND2_X1 U539 ( .A1(n420), .A2(n604), .ZN(n419) );
  NAND2_X1 U540 ( .A1(n422), .A2(n535), .ZN(n421) );
  NAND2_X1 U541 ( .A1(n427), .A2(n426), .ZN(n422) );
  NAND2_X1 U542 ( .A1(n650), .A2(n430), .ZN(n427) );
  NOR2_X1 U543 ( .A1(n650), .A2(KEYINPUT75), .ZN(n534) );
  INV_X1 U544 ( .A(KEYINPUT75), .ZN(n429) );
  XNOR2_X2 U545 ( .A(n507), .B(n506), .ZN(n431) );
  NOR2_X2 U546 ( .A1(n634), .A2(n755), .ZN(n597) );
  NAND2_X1 U547 ( .A1(n436), .A2(n435), .ZN(n434) );
  AND2_X1 U548 ( .A1(n599), .A2(n437), .ZN(n634) );
  NOR2_X1 U549 ( .A1(n591), .A2(n600), .ZN(n437) );
  NOR2_X1 U550 ( .A1(n592), .A2(n590), .ZN(n599) );
  INV_X1 U551 ( .A(KEYINPUT12), .ZN(n511) );
  INV_X1 U552 ( .A(KEYINPUT36), .ZN(n543) );
  INV_X1 U553 ( .A(n612), .ZN(n613) );
  INV_X1 U554 ( .A(KEYINPUT41), .ZN(n561) );
  XNOR2_X1 U555 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U556 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U557 ( .A(n724), .B(n723), .ZN(n725) );
  XOR2_X1 U558 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n439) );
  NAND2_X1 U559 ( .A1(G234), .A2(n612), .ZN(n438) );
  XNOR2_X1 U560 ( .A(n439), .B(n438), .ZN(n459) );
  NAND2_X1 U561 ( .A1(n459), .A2(G221), .ZN(n440) );
  XOR2_X1 U562 ( .A(KEYINPUT21), .B(n440), .Z(n441) );
  XNOR2_X1 U563 ( .A(KEYINPUT92), .B(n441), .ZN(n678) );
  XNOR2_X1 U564 ( .A(n442), .B(KEYINPUT14), .ZN(n445) );
  NAND2_X1 U565 ( .A1(G902), .A2(n445), .ZN(n578) );
  NOR2_X1 U566 ( .A1(G900), .A2(n578), .ZN(n443) );
  NAND2_X1 U567 ( .A1(G953), .A2(n443), .ZN(n444) );
  XNOR2_X1 U568 ( .A(n444), .B(KEYINPUT101), .ZN(n446) );
  NAND2_X1 U569 ( .A1(G952), .A2(n445), .ZN(n701) );
  NOR2_X1 U570 ( .A1(n701), .A2(G953), .ZN(n580) );
  NOR2_X1 U571 ( .A1(n446), .A2(n580), .ZN(n548) );
  INV_X2 U572 ( .A(G953), .ZN(n746) );
  NAND2_X1 U573 ( .A1(n524), .A2(G221), .ZN(n448) );
  XOR2_X1 U574 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n450) );
  XNOR2_X1 U575 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U576 ( .A(n744), .B(n451), .ZN(n452) );
  XNOR2_X1 U577 ( .A(n453), .B(n452), .ZN(n456) );
  XOR2_X1 U578 ( .A(G119), .B(G110), .Z(n734) );
  INV_X1 U579 ( .A(n734), .ZN(n454) );
  XNOR2_X1 U580 ( .A(G137), .B(n497), .ZN(n455) );
  XNOR2_X1 U581 ( .A(n456), .B(n455), .ZN(n722) );
  INV_X1 U582 ( .A(n722), .ZN(n458) );
  NAND2_X1 U583 ( .A1(n459), .A2(G217), .ZN(n461) );
  XNOR2_X1 U584 ( .A(KEYINPUT25), .B(KEYINPUT79), .ZN(n460) );
  XNOR2_X2 U585 ( .A(n463), .B(n462), .ZN(n600) );
  XNOR2_X1 U586 ( .A(n492), .B(n466), .ZN(n467) );
  XNOR2_X1 U587 ( .A(n470), .B(n469), .ZN(n474) );
  NOR2_X2 U588 ( .A1(G953), .A2(G237), .ZN(n508) );
  NAND2_X1 U589 ( .A1(G210), .A2(n508), .ZN(n472) );
  XNOR2_X1 U590 ( .A(n473), .B(n474), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n488), .B(n475), .ZN(n476) );
  INV_X1 U592 ( .A(n476), .ZN(n477) );
  INV_X1 U593 ( .A(KEYINPUT28), .ZN(n478) );
  NAND2_X1 U594 ( .A1(G227), .A2(n746), .ZN(n480) );
  XNOR2_X1 U595 ( .A(n487), .B(n481), .ZN(n482) );
  XNOR2_X1 U596 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n743), .B(n484), .ZN(n624) );
  NAND2_X1 U598 ( .A1(n624), .A2(n457), .ZN(n486) );
  XOR2_X1 U599 ( .A(KEYINPUT70), .B(G469), .Z(n485) );
  XOR2_X1 U600 ( .A(KEYINPUT17), .B(G125), .Z(n494) );
  NAND2_X1 U601 ( .A1(G224), .A2(n746), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n496), .B(KEYINPUT18), .ZN(n498) );
  NAND2_X1 U603 ( .A1(n636), .A2(n612), .ZN(n501) );
  NAND2_X1 U604 ( .A1(n457), .A2(n499), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n502), .A2(G210), .ZN(n500) );
  INV_X1 U606 ( .A(n557), .ZN(n503) );
  NAND2_X1 U607 ( .A1(n502), .A2(G214), .ZN(n670) );
  NAND2_X1 U608 ( .A1(n503), .A2(n670), .ZN(n507) );
  XOR2_X1 U609 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n505) );
  INV_X1 U610 ( .A(KEYINPUT19), .ZN(n504) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(G475), .ZN(n522) );
  NAND2_X1 U612 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n513) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n515) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U616 ( .A(n744), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U618 ( .A(n520), .B(n519), .ZN(n712) );
  NOR2_X1 U619 ( .A1(G902), .A2(n712), .ZN(n521) );
  XNOR2_X1 U620 ( .A(n522), .B(n521), .ZN(n559) );
  INV_X1 U621 ( .A(KEYINPUT98), .ZN(n523) );
  XNOR2_X1 U622 ( .A(n559), .B(n523), .ZN(n532) );
  NAND2_X1 U623 ( .A1(G217), .A2(n524), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n529), .B(n530), .ZN(n718) );
  NAND2_X1 U626 ( .A1(n718), .A2(n457), .ZN(n531) );
  INV_X1 U627 ( .A(n660), .ZN(n533) );
  NAND2_X1 U628 ( .A1(KEYINPUT47), .A2(n534), .ZN(n536) );
  INV_X1 U629 ( .A(KEYINPUT81), .ZN(n535) );
  NOR2_X1 U630 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U631 ( .A(n538), .ZN(n569) );
  BUF_X1 U632 ( .A(n557), .Z(n539) );
  INV_X1 U633 ( .A(n654), .ZN(n657) );
  XNOR2_X1 U634 ( .A(n683), .B(KEYINPUT6), .ZN(n598) );
  NAND2_X1 U635 ( .A1(n542), .A2(n670), .ZN(n571) );
  XNOR2_X2 U636 ( .A(n549), .B(KEYINPUT1), .ZN(n686) );
  XNOR2_X1 U637 ( .A(n686), .B(KEYINPUT86), .ZN(n593) );
  NOR2_X1 U638 ( .A1(n546), .A2(n593), .ZN(n664) );
  NAND2_X1 U639 ( .A1(KEYINPUT81), .A2(n674), .ZN(n547) );
  NOR2_X1 U640 ( .A1(n687), .A2(n548), .ZN(n550) );
  INV_X1 U641 ( .A(n549), .ZN(n604) );
  NAND2_X1 U642 ( .A1(n550), .A2(n604), .ZN(n553) );
  XNOR2_X1 U643 ( .A(n551), .B(KEYINPUT30), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n586) );
  NOR2_X1 U645 ( .A1(n539), .A2(n586), .ZN(n554) );
  NAND2_X1 U646 ( .A1(n565), .A2(n554), .ZN(n630) );
  XOR2_X1 U647 ( .A(KEYINPUT82), .B(n630), .Z(n555) );
  XNOR2_X1 U648 ( .A(n557), .B(KEYINPUT38), .ZN(n669) );
  NAND2_X1 U649 ( .A1(n670), .A2(n669), .ZN(n558) );
  NOR2_X1 U650 ( .A1(n560), .A2(n559), .ZN(n671) );
  NAND2_X1 U651 ( .A1(n673), .A2(n671), .ZN(n562) );
  XOR2_X1 U652 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n566) );
  XOR2_X1 U653 ( .A(KEYINPUT69), .B(KEYINPUT48), .Z(n570) );
  INV_X1 U654 ( .A(n686), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n572), .B(KEYINPUT43), .ZN(n573) );
  AND2_X1 U656 ( .A1(n539), .A2(n573), .ZN(n574) );
  INV_X1 U657 ( .A(n575), .ZN(n576) );
  NOR2_X1 U658 ( .A1(n576), .A2(n660), .ZN(n631) );
  XNOR2_X1 U659 ( .A(KEYINPUT87), .B(G898), .ZN(n730) );
  NAND2_X1 U660 ( .A1(n730), .A2(G953), .ZN(n577) );
  XNOR2_X1 U661 ( .A(n577), .B(KEYINPUT88), .ZN(n738) );
  NOR2_X1 U662 ( .A1(n578), .A2(n738), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X2 U664 ( .A(n582), .B(KEYINPUT0), .ZN(n607) );
  INV_X1 U665 ( .A(n602), .ZN(n583) );
  NOR2_X1 U666 ( .A1(n583), .A2(n598), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n584), .B(KEYINPUT33), .ZN(n703) );
  INV_X1 U668 ( .A(n600), .ZN(n679) );
  NAND2_X1 U669 ( .A1(n671), .A2(n678), .ZN(n587) );
  NOR2_X1 U670 ( .A1(n592), .A2(n600), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n593), .A2(n375), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X2 U673 ( .A(n596), .B(KEYINPUT32), .ZN(n758) );
  AND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n643) );
  NAND2_X1 U676 ( .A1(n602), .A2(n683), .ZN(n692) );
  NOR2_X1 U677 ( .A1(n607), .A2(n692), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT31), .B(n603), .ZN(n659) );
  NOR2_X1 U679 ( .A1(n687), .A2(n683), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  OR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n646) );
  NAND2_X1 U682 ( .A1(n659), .A2(n646), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n608), .A2(n674), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n727) );
  XNOR2_X1 U686 ( .A(n666), .B(KEYINPUT2), .ZN(n614) );
  AND2_X2 U687 ( .A1(n614), .A2(n613), .ZN(n720) );
  NAND2_X1 U688 ( .A1(n720), .A2(G472), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT62), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(n619) );
  INV_X1 U691 ( .A(G952), .ZN(n618) );
  NOR2_X2 U692 ( .A1(n619), .A2(n726), .ZN(n621) );
  XNOR2_X1 U693 ( .A(KEYINPUT63), .B(KEYINPUT85), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(G57) );
  NAND2_X1 U695 ( .A1(n720), .A2(G469), .ZN(n626) );
  XNOR2_X1 U696 ( .A(KEYINPUT58), .B(KEYINPUT116), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT57), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U700 ( .A1(n627), .A2(n726), .ZN(n629) );
  INV_X1 U701 ( .A(KEYINPUT117), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(G54) );
  XNOR2_X1 U703 ( .A(n630), .B(G143), .ZN(G45) );
  XOR2_X1 U704 ( .A(G134), .B(n631), .Z(G36) );
  XOR2_X1 U705 ( .A(G131), .B(KEYINPUT126), .Z(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(G33) );
  XOR2_X1 U707 ( .A(G110), .B(n634), .Z(G12) );
  NAND2_X1 U708 ( .A1(n720), .A2(G210), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(n640) );
  INV_X1 U712 ( .A(n726), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n642) );
  INV_X1 U714 ( .A(KEYINPUT56), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G51) );
  XNOR2_X1 U716 ( .A(G101), .B(n643), .ZN(G3) );
  NOR2_X1 U717 ( .A1(n657), .A2(n646), .ZN(n645) );
  XNOR2_X1 U718 ( .A(G104), .B(KEYINPUT107), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(G6) );
  NOR2_X1 U720 ( .A1(n660), .A2(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U723 ( .A(G107), .B(n649), .ZN(G9) );
  NOR2_X1 U724 ( .A1(n660), .A2(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(KEYINPUT29), .B(KEYINPUT108), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(G128), .B(n653), .ZN(G30) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(G146), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n657), .A2(n659), .ZN(n658) );
  XOR2_X1 U731 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n662) );
  XNOR2_X1 U733 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(G116), .B(n663), .ZN(G18) );
  XNOR2_X1 U736 ( .A(G125), .B(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U738 ( .A1(n666), .A2(KEYINPUT80), .ZN(n668) );
  INV_X1 U739 ( .A(KEYINPUT2), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n708) );
  OR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n677), .A2(n703), .ZN(n698) );
  INV_X1 U746 ( .A(n678), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT49), .ZN(n682) );
  XNOR2_X1 U749 ( .A(KEYINPUT111), .B(n682), .ZN(n685) );
  INV_X1 U750 ( .A(n683), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n690) );
  NAND2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U753 ( .A(KEYINPUT50), .B(n688), .Z(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U755 ( .A(KEYINPUT112), .B(n691), .Z(n693) );
  NAND2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n695) );
  XOR2_X1 U757 ( .A(KEYINPUT51), .B(KEYINPUT113), .Z(n694) );
  XNOR2_X1 U758 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n696), .A2(n702), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT52), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U765 ( .A(KEYINPUT114), .B(n706), .Z(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n709), .B(KEYINPUT115), .ZN(n710) );
  NOR2_X1 U768 ( .A1(G953), .A2(n710), .ZN(n711) );
  XNOR2_X1 U769 ( .A(KEYINPUT53), .B(n711), .ZN(G75) );
  NAND2_X1 U770 ( .A1(n720), .A2(G475), .ZN(n714) );
  XOR2_X1 U771 ( .A(n712), .B(KEYINPUT59), .Z(n713) );
  XNOR2_X1 U772 ( .A(n716), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U773 ( .A1(n720), .A2(G478), .ZN(n717) );
  XOR2_X1 U774 ( .A(n718), .B(n717), .Z(n719) );
  NOR2_X1 U775 ( .A1(n726), .A2(n719), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n720), .A2(G217), .ZN(n724) );
  XOR2_X1 U777 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n721) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(G66) );
  XNOR2_X1 U779 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n742) );
  NAND2_X1 U780 ( .A1(n727), .A2(n746), .ZN(n733) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(n728), .Z(n729) );
  NOR2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U784 ( .A(KEYINPUT120), .B(n731), .Z(n732) );
  NAND2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n740) );
  XOR2_X1 U786 ( .A(n735), .B(n356), .Z(n736) );
  XNOR2_X1 U787 ( .A(KEYINPUT121), .B(n736), .ZN(n737) );
  NAND2_X1 U788 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(G69) );
  XOR2_X1 U791 ( .A(n743), .B(n744), .Z(n749) );
  XNOR2_X1 U792 ( .A(n745), .B(n749), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U794 ( .A(n748), .B(KEYINPUT124), .ZN(n753) );
  XOR2_X1 U795 ( .A(G227), .B(n749), .Z(n750) );
  NAND2_X1 U796 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U797 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(n754), .Z(G72) );
  XOR2_X1 U800 ( .A(n755), .B(G122), .Z(G24) );
  XOR2_X1 U801 ( .A(n756), .B(G137), .Z(G39) );
  XOR2_X1 U802 ( .A(G140), .B(n757), .Z(G42) );
  XNOR2_X1 U803 ( .A(n758), .B(G119), .ZN(G21) );
endmodule

