

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X2 U323 ( .A(n473), .B(KEYINPUT99), .ZN(n483) );
  NOR2_X2 U324 ( .A1(n500), .A2(n567), .ZN(n497) );
  XNOR2_X1 U325 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U326 ( .A(n318), .B(n317), .ZN(n356) );
  INV_X1 U327 ( .A(n467), .ZN(n468) );
  XNOR2_X1 U328 ( .A(n466), .B(KEYINPUT97), .ZN(n469) );
  NAND2_X1 U329 ( .A1(n475), .A2(n582), .ZN(n476) );
  XNOR2_X1 U330 ( .A(n474), .B(KEYINPUT103), .ZN(n475) );
  XOR2_X1 U331 ( .A(n409), .B(n408), .Z(n463) );
  XNOR2_X1 U332 ( .A(n352), .B(n351), .ZN(n355) );
  XNOR2_X1 U333 ( .A(n326), .B(n325), .ZN(n519) );
  NOR2_X1 U334 ( .A1(n463), .A2(n429), .ZN(n291) );
  XOR2_X1 U335 ( .A(n299), .B(n298), .Z(n292) );
  INV_X1 U336 ( .A(KEYINPUT84), .ZN(n396) );
  XNOR2_X1 U337 ( .A(n397), .B(n396), .ZN(n398) );
  AND2_X1 U338 ( .A1(n469), .A2(n468), .ZN(n470) );
  INV_X1 U339 ( .A(G64GAT), .ZN(n315) );
  XNOR2_X1 U340 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U341 ( .A(n316), .B(n315), .ZN(n318) );
  XNOR2_X1 U342 ( .A(n387), .B(KEYINPUT121), .ZN(n388) );
  XNOR2_X1 U343 ( .A(n300), .B(n292), .ZN(n301) );
  XNOR2_X1 U344 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n377) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U346 ( .A(KEYINPUT36), .B(n555), .Z(n582) );
  XNOR2_X1 U347 ( .A(n575), .B(n377), .ZN(n503) );
  XNOR2_X1 U348 ( .A(n476), .B(KEYINPUT37), .ZN(n516) );
  XNOR2_X1 U349 ( .A(KEYINPUT91), .B(n467), .ZN(n567) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n555) );
  INV_X1 U351 ( .A(G43GAT), .ZN(n478) );
  XNOR2_X1 U352 ( .A(n447), .B(G190GAT), .ZN(n448) );
  XNOR2_X1 U353 ( .A(n478), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U354 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XNOR2_X1 U355 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U356 ( .A(G85GAT), .B(G99GAT), .Z(n344) );
  XOR2_X1 U357 ( .A(G190GAT), .B(G36GAT), .Z(n319) );
  XOR2_X1 U358 ( .A(n344), .B(n319), .Z(n294) );
  NAND2_X1 U359 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U360 ( .A(n294), .B(n293), .ZN(n302) );
  XOR2_X1 U361 ( .A(G29GAT), .B(G134GAT), .Z(n418) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G106GAT), .Z(n296) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U364 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U365 ( .A(n418), .B(n297), .ZN(n300) );
  XOR2_X1 U366 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n299) );
  XNOR2_X1 U367 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n298) );
  XOR2_X1 U368 ( .A(n303), .B(KEYINPUT10), .Z(n307) );
  XOR2_X1 U369 ( .A(G43GAT), .B(G50GAT), .Z(n305) );
  XNOR2_X1 U370 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n304) );
  XNOR2_X1 U371 ( .A(n305), .B(n304), .ZN(n371) );
  XNOR2_X1 U372 ( .A(n371), .B(KEYINPUT9), .ZN(n306) );
  XOR2_X1 U373 ( .A(G169GAT), .B(KEYINPUT19), .Z(n309) );
  XNOR2_X1 U374 ( .A(G183GAT), .B(KEYINPUT81), .ZN(n308) );
  XNOR2_X1 U375 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U376 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n310) );
  XOR2_X1 U377 ( .A(n311), .B(n310), .Z(n443) );
  XOR2_X1 U378 ( .A(KEYINPUT21), .B(G197GAT), .Z(n313) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(KEYINPUT85), .ZN(n312) );
  XNOR2_X1 U380 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U381 ( .A(G211GAT), .B(n314), .Z(n401) );
  XNOR2_X1 U382 ( .A(n443), .B(n401), .ZN(n326) );
  XNOR2_X1 U383 ( .A(G92GAT), .B(G176GAT), .ZN(n316) );
  XOR2_X1 U384 ( .A(G204GAT), .B(KEYINPUT72), .Z(n317) );
  XOR2_X1 U385 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n321) );
  XNOR2_X1 U386 ( .A(n319), .B(G8GAT), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U388 ( .A(n356), .B(n322), .Z(n324) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G15GAT), .Z(n328) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n370) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n329), .B(KEYINPUT69), .ZN(n357) );
  XNOR2_X1 U396 ( .A(n370), .B(n357), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n331) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U400 ( .A(n332), .B(KEYINPUT12), .Z(n340) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G211GAT), .Z(n334) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U403 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U404 ( .A(KEYINPUT14), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U405 ( .A(G57GAT), .B(G183GAT), .ZN(n335) );
  XNOR2_X1 U406 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U407 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U409 ( .A(n342), .B(n341), .Z(n579) );
  NAND2_X1 U410 ( .A1(n582), .A2(n579), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n343), .B(KEYINPUT45), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n346) );
  XOR2_X1 U413 ( .A(G120GAT), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U414 ( .A(n413), .B(n344), .ZN(n345) );
  XNOR2_X1 U415 ( .A(n346), .B(n345), .ZN(n352) );
  XOR2_X1 U416 ( .A(KEYINPUT71), .B(KEYINPUT74), .Z(n348) );
  XNOR2_X1 U417 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n347) );
  XNOR2_X1 U418 ( .A(n348), .B(n347), .ZN(n350) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XOR2_X1 U420 ( .A(KEYINPUT70), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U421 ( .A(G148GAT), .B(G106GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n399) );
  XNOR2_X1 U423 ( .A(n355), .B(n399), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n575) );
  NOR2_X1 U426 ( .A1(n360), .A2(n575), .ZN(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT114), .B(n361), .ZN(n376) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G29GAT), .Z(n363) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n365) );
  XNOR2_X1 U432 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U434 ( .A(G197GAT), .B(G169GAT), .Z(n367) );
  XNOR2_X1 U435 ( .A(G141GAT), .B(G113GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U437 ( .A(n369), .B(n368), .Z(n373) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n571) );
  INV_X1 U441 ( .A(n571), .ZN(n544) );
  NAND2_X1 U442 ( .A1(n376), .A2(n544), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n544), .A2(n503), .ZN(n379) );
  INV_X1 U444 ( .A(KEYINPUT46), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  INV_X1 U446 ( .A(n579), .ZN(n565) );
  NAND2_X1 U447 ( .A1(n380), .A2(n565), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n381), .B(KEYINPUT113), .ZN(n382) );
  NAND2_X1 U449 ( .A1(n382), .A2(n555), .ZN(n383) );
  XOR2_X1 U450 ( .A(KEYINPUT47), .B(n383), .Z(n384) );
  NAND2_X1 U451 ( .A1(n385), .A2(n384), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT48), .B(n386), .Z(n528) );
  NOR2_X1 U453 ( .A1(n519), .A2(n528), .ZN(n389) );
  INV_X1 U454 ( .A(KEYINPUT54), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n568) );
  XOR2_X1 U456 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n391) );
  XNOR2_X1 U457 ( .A(G50GAT), .B(G22GAT), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U459 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n393) );
  XNOR2_X1 U460 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U462 ( .A(n395), .B(n394), .Z(n403) );
  NAND2_X1 U463 ( .A1(G228GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n409) );
  XNOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n404), .B(KEYINPUT3), .ZN(n405) );
  XOR2_X1 U468 ( .A(n405), .B(KEYINPUT86), .Z(n407) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(G162GAT), .ZN(n406) );
  XOR2_X1 U470 ( .A(n407), .B(n406), .Z(n426) );
  INV_X1 U471 ( .A(n426), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n411) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U475 ( .A(n412), .B(G148GAT), .Z(n415) );
  XNOR2_X1 U476 ( .A(n413), .B(G85GAT), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n422) );
  XOR2_X1 U478 ( .A(G113GAT), .B(G127GAT), .Z(n417) );
  XNOR2_X1 U479 ( .A(KEYINPUT80), .B(KEYINPUT0), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n440) );
  XOR2_X1 U481 ( .A(n418), .B(n440), .Z(n420) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n424) );
  XNOR2_X1 U486 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U488 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n467) );
  INV_X1 U490 ( .A(n567), .ZN(n429) );
  AND2_X1 U491 ( .A1(n568), .A2(n291), .ZN(n430) );
  XOR2_X1 U492 ( .A(KEYINPUT55), .B(n430), .Z(n446) );
  XOR2_X1 U493 ( .A(G43GAT), .B(G134GAT), .Z(n432) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U496 ( .A(G176GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G120GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U499 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U500 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n438) );
  XNOR2_X1 U501 ( .A(G99GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X2 U505 ( .A(n444), .B(n443), .Z(n531) );
  INV_X1 U506 ( .A(n531), .ZN(n445) );
  NAND2_X1 U507 ( .A1(n446), .A2(n445), .ZN(n564) );
  NOR2_X1 U508 ( .A1(n555), .A2(n564), .ZN(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n447) );
  NOR2_X1 U510 ( .A1(n544), .A2(n564), .ZN(n452) );
  INV_X1 U511 ( .A(KEYINPUT122), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n450), .B(G169GAT), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(G1348GAT) );
  NOR2_X1 U514 ( .A1(n544), .A2(n575), .ZN(n453) );
  XOR2_X1 U515 ( .A(KEYINPUT75), .B(n453), .Z(n486) );
  XNOR2_X1 U516 ( .A(n519), .B(KEYINPUT27), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n454), .B(KEYINPUT94), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n463), .B(KEYINPUT28), .ZN(n455) );
  XOR2_X2 U519 ( .A(n455), .B(KEYINPUT66), .Z(n525) );
  INV_X1 U520 ( .A(n525), .ZN(n456) );
  NOR2_X1 U521 ( .A1(n461), .A2(n456), .ZN(n529) );
  NAND2_X1 U522 ( .A1(n531), .A2(n529), .ZN(n457) );
  NOR2_X1 U523 ( .A1(n567), .A2(n457), .ZN(n458) );
  XOR2_X1 U524 ( .A(KEYINPUT95), .B(n458), .Z(n472) );
  NAND2_X1 U525 ( .A1(n463), .A2(n531), .ZN(n459) );
  XNOR2_X1 U526 ( .A(n459), .B(KEYINPUT26), .ZN(n460) );
  XNOR2_X1 U527 ( .A(KEYINPUT96), .B(n460), .ZN(n570) );
  NOR2_X1 U528 ( .A1(n461), .A2(n570), .ZN(n543) );
  NOR2_X1 U529 ( .A1(n531), .A2(n519), .ZN(n462) );
  NOR2_X1 U530 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NOR2_X1 U532 ( .A1(n543), .A2(n465), .ZN(n466) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(n470), .ZN(n471) );
  NOR2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n483), .A2(n565), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n486), .A2(n516), .ZN(n477) );
  XNOR2_X2 U537 ( .A(n477), .B(KEYINPUT38), .ZN(n500) );
  NOR2_X1 U538 ( .A1(n531), .A2(n500), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n579), .A2(n555), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT16), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT79), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(n485), .Z(n504) );
  NAND2_X1 U544 ( .A1(n486), .A2(n504), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n567), .A2(n494), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n519), .A2(n494), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT102), .B(n490), .Z(n491) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U552 ( .A1(n531), .A2(n494), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n525), .A2(n494), .ZN(n495) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n519), .A2(n500), .ZN(n499) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n500), .A2(n525), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT106), .ZN(n558) );
  NOR2_X1 U566 ( .A1(n571), .A2(n558), .ZN(n515) );
  NAND2_X1 U567 ( .A1(n515), .A2(n504), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n567), .A2(n511), .ZN(n505) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n511), .ZN(n507) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n531), .A2(n511), .ZN(n508) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n510) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(n513) );
  NOR2_X1 U578 ( .A1(n525), .A2(n511), .ZN(n512) );
  XOR2_X1 U579 ( .A(n513), .B(n512), .Z(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT107), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n567), .A2(n524), .ZN(n517) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n517), .Z(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT110), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n524), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n531), .A2(n524), .ZN(n523) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n567), .A2(n528), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n529), .A2(n542), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n535), .A2(n571), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  INV_X1 U599 ( .A(n535), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n558), .A2(n539), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U604 ( .A1(n535), .A2(n579), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n555), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n544), .A2(n554), .ZN(n545) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n503), .A2(n554), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(KEYINPUT52), .B(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n565), .A2(n554), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n564), .A2(n558), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n560) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n583), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n583), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

