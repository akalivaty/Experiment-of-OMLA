//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT28), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR3_X1   g008(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT70), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT27), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n212), .B1(new_n215), .B2(new_n203), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G190gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT27), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n209), .B1(new_n221), .B2(new_n215), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n210), .A2(new_n218), .B1(new_n222), .B2(KEYINPUT28), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT71), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n220), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n205), .B1(new_n229), .B2(KEYINPUT27), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n212), .B1(new_n230), .B2(new_n209), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT70), .B1(new_n206), .B2(new_n209), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n211), .A3(new_n217), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n234), .A3(KEYINPUT71), .ZN(new_n235));
  INV_X1    g034(.A(G169gat), .ZN(new_n236));
  INV_X1    g035(.A(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239));
  OR3_X1    g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT26), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n238), .B2(KEYINPUT26), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(KEYINPUT26), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n225), .A2(new_n226), .A3(new_n235), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n248), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n250), .B(new_n252), .C1(new_n209), .C2(new_n229), .ZN(new_n253));
  OR2_X1    g052(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n238), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT23), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n256), .A2(new_n243), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n258), .A3(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n257), .B(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n252), .B(new_n246), .C1(G183gat), .C2(G190gat), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n262), .A2(new_n243), .A3(new_n256), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n253), .A2(new_n258), .A3(new_n267), .A4(KEYINPUT25), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n245), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n272), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n245), .A2(new_n276), .A3(new_n269), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G227gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n202), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n278), .A2(KEYINPUT34), .A3(new_n285), .A4(new_n279), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(KEYINPUT75), .A3(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n245), .A2(new_n276), .A3(new_n269), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n276), .B1(new_n245), .B2(new_n269), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(KEYINPUT32), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G15gat), .B(G43gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n280), .B2(new_n283), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(KEYINPUT33), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND4_X1   g100(.A1(new_n297), .A2(new_n290), .A3(KEYINPUT32), .A4(new_n300), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n287), .B(new_n296), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT75), .B1(new_n284), .B2(new_n286), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n297), .A3(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n304), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n287), .A4(new_n296), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(G141gat), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT2), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G155gat), .B(G162gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT80), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n320), .A2(new_n327), .A3(new_n323), .A4(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n318), .A2(G148gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT2), .B1(new_n317), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(new_n324), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT81), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  AOI211_X1 g134(.A(new_n335), .B(new_n332), .C1(new_n326), .C2(new_n328), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n277), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n326), .B2(new_n328), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n276), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT82), .Z(new_n342));
  AOI21_X1  g141(.A(new_n313), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(new_n334), .B2(new_n336), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n277), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n339), .B(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(new_n338), .B2(new_n276), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n343), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n347), .A2(new_n348), .A3(new_n313), .A4(new_n350), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n362), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n358), .B1(new_n352), .B2(new_n353), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT83), .B1(new_n366), .B2(KEYINPUT6), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  INV_X1    g170(.A(G92gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT76), .B(G64gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  XOR2_X1   g174(.A(G197gat), .B(G204gat), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G211gat), .A2(G218gat), .ZN(new_n378));
  OR2_X1    g177(.A1(G211gat), .A2(G218gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n378), .B(new_n379), .C1(new_n376), .C2(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT29), .B(new_n387), .C1(new_n245), .C2(new_n269), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n245), .A2(new_n387), .A3(new_n269), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n270), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n245), .A2(new_n387), .A3(new_n269), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n384), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n375), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n370), .B1(new_n395), .B2(KEYINPUT30), .ZN(new_n396));
  INV_X1    g195(.A(new_n375), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n388), .A2(new_n385), .A3(new_n389), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n384), .B1(new_n392), .B2(new_n393), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT78), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n398), .A2(new_n399), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n375), .B(KEYINPUT77), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n400), .B2(new_n401), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n383), .B(KEYINPUT85), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n382), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n411), .B2(new_n391), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n412), .B2(new_n338), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n384), .B1(new_n346), .B2(new_n391), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n334), .A2(new_n336), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT3), .B1(new_n384), .B2(new_n391), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n414), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n413), .A2(new_n414), .B1(new_n418), .B2(new_n409), .ZN(new_n419));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G22gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422));
  INV_X1    g221(.A(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n421), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n419), .B(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n312), .A2(new_n369), .A3(new_n408), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT35), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n427), .B2(KEYINPUT35), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n352), .A2(KEYINPUT87), .A3(new_n353), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT87), .B1(new_n352), .B2(new_n353), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n359), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n365), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n433), .A2(new_n434), .B1(KEYINPUT6), .B2(new_n366), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n403), .B2(new_n407), .ZN(new_n438));
  AOI22_X1  g237(.A1(KEYINPUT30), .A2(new_n395), .B1(new_n404), .B2(new_n405), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT86), .A3(new_n396), .A4(new_n402), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n426), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n305), .B2(new_n311), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n436), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n429), .A2(new_n430), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n354), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n352), .A2(KEYINPUT87), .A3(new_n353), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n350), .B1(new_n347), .B2(new_n348), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n340), .A2(new_n342), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(KEYINPUT39), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n358), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n358), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n450), .A2(new_n456), .A3(new_n452), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT40), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n449), .A2(new_n359), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n440), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT88), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n390), .A2(KEYINPUT37), .A3(new_n394), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n375), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n390), .B2(new_n394), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT38), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n405), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n465), .B(new_n471), .C1(new_n404), .C2(new_n467), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n469), .A2(new_n400), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n442), .B1(new_n435), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n438), .A2(new_n462), .A3(new_n475), .A4(new_n440), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n464), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n426), .B1(new_n369), .B2(new_n408), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n311), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT36), .B1(new_n305), .B2(new_n311), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n445), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT8), .ZN(new_n486));
  NAND2_X1  g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G85gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n372), .ZN(new_n491));
  NAND3_X1  g290(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n492));
  AND4_X1   g291(.A1(new_n486), .A2(new_n489), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT104), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G99gat), .ZN(new_n497));
  INV_X1    g296(.A(G106gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT104), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n485), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT105), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n493), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n493), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT106), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n493), .A2(new_n502), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT105), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT106), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n502), .A3(new_n503), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n493), .A2(new_n502), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT100), .B(G57gat), .ZN(new_n514));
  INV_X1    g313(.A(G64gat), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT101), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G57gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(G64gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT101), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n517), .A2(KEYINPUT100), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n517), .A2(KEYINPUT100), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n520), .B(G64gat), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT102), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT9), .ZN(new_n527));
  INV_X1    g326(.A(G71gat), .ZN(new_n528));
  INV_X1    g327(.A(G78gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n525), .B(KEYINPUT99), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n515), .A2(G57gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT10), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n508), .A2(new_n510), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n512), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT103), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n531), .A2(KEYINPUT103), .A3(new_n535), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT10), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n542), .A2(new_n548), .B1(G230gat), .B2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n537), .B2(new_n541), .ZN(new_n551));
  XNOR2_X1  g350(.A(G120gat), .B(G148gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G176gat), .B(G204gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n549), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n550), .B(KEYINPUT107), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n542), .B2(new_n548), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n554), .B1(new_n559), .B2(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n484), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n544), .B2(new_n545), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(G1gat), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n569), .A2(G183gat), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(G183gat), .B1(new_n569), .B2(new_n578), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n567), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n581), .A3(new_n567), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(G231gat), .A4(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n584), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n582), .ZN(new_n588));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G211gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n585), .B2(new_n588), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n565), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n564), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G29gat), .A2(G36gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT92), .ZN(new_n600));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT15), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT14), .ZN(new_n606));
  INV_X1    g405(.A(G29gat), .ZN(new_n607));
  INV_X1    g406(.A(G36gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT15), .B1(new_n601), .B2(KEYINPUT94), .ZN(new_n612));
  AND4_X1   g411(.A1(new_n600), .A2(new_n605), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n610), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(G29gat), .A2(G36gat), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT91), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n600), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n604), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT93), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n622), .A3(new_n619), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n613), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n577), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n612), .A3(new_n600), .A4(new_n611), .ZN(new_n626));
  INV_X1    g425(.A(new_n623), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n578), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n630), .A3(KEYINPUT96), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n624), .A2(KEYINPUT96), .A3(new_n577), .ZN(new_n632));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n631), .A2(new_n632), .A3(new_n638), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT11), .B(G169gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  INV_X1    g445(.A(new_n630), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT17), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n624), .B2(KEYINPUT95), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n629), .A2(new_n650), .A3(KEYINPUT17), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n652), .B2(new_n577), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n646), .B1(new_n653), .B2(new_n633), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n578), .B1(new_n649), .B2(new_n651), .ZN(new_n655));
  INV_X1    g454(.A(new_n633), .ZN(new_n656));
  NOR4_X1   g455(.A1(new_n655), .A2(KEYINPUT18), .A3(new_n656), .A4(new_n647), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n640), .B(new_n645), .C1(new_n654), .C2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n652), .A2(new_n577), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n633), .A3(new_n630), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT18), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n646), .A3(new_n633), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n645), .A4(new_n640), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n640), .ZN(new_n668));
  INV_X1    g467(.A(new_n645), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n513), .ZN(new_n673));
  NAND3_X1  g472(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n547), .A2(new_n629), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G190gat), .B(G218gat), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(G134gat), .B(G162gat), .Z(new_n679));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n678), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n598), .A2(new_n672), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n563), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n369), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  INV_X1    g490(.A(new_n441), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n573), .A2(new_n572), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n563), .A2(new_n686), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n573), .A2(new_n572), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G8gat), .B1(new_n687), .B2(new_n441), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(G1325gat));
  NOR2_X1   g499(.A1(new_n480), .A2(new_n481), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n688), .A2(G15gat), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n688), .B2(new_n312), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n426), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n598), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n672), .A3(new_n561), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n484), .A2(new_n685), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n607), .A3(new_n689), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n685), .B1(new_n445), .B2(new_n483), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT44), .B(new_n685), .C1(new_n445), .C2(new_n483), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n720), .A2(new_n689), .A3(new_n710), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n713), .B1(new_n607), .B2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n711), .A2(new_n608), .A3(new_n692), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT46), .Z(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n692), .A3(new_n710), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G36gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1329gat));
  NAND4_X1  g526(.A1(new_n716), .A2(new_n702), .A3(new_n718), .A4(new_n710), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  INV_X1    g528(.A(G43gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n730), .A3(new_n312), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1330gat));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n442), .A3(new_n718), .A4(new_n710), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G50gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n423), .A3(new_n442), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1331gat));
  INV_X1    g539(.A(new_n685), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n709), .A2(new_n672), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n484), .A2(new_n561), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n369), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(new_n514), .Z(G1332gat));
  OR2_X1    g545(.A1(new_n744), .A2(new_n441), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  OAI21_X1  g550(.A(G71gat), .B1(new_n744), .B2(new_n701), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n312), .A2(new_n528), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n484), .A2(new_n561), .A3(new_n743), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n752), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n752), .A2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(KEYINPUT50), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1334gat));
  NOR2_X1   g563(.A1(new_n744), .A2(new_n426), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n529), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n709), .A2(new_n671), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n685), .B(new_n767), .C1(new_n445), .C2(new_n483), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(KEYINPUT51), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n561), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n771), .A2(new_n369), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n561), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n717), .A2(new_n719), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n369), .A2(new_n490), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n772), .A2(new_n490), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  INV_X1    g575(.A(new_n773), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n716), .A2(new_n692), .A3(new_n718), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n692), .A2(new_n372), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n779), .B(new_n780), .C1(new_n771), .C2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n778), .A2(new_n783), .A3(G92gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n778), .B2(G92gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n441), .A2(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n561), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n768), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n788), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n784), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n782), .B1(new_n792), .B2(new_n780), .ZN(G1337gat));
  NAND4_X1  g592(.A1(new_n716), .A2(new_n702), .A3(new_n718), .A4(new_n777), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(G99gat), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n312), .A2(new_n497), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n771), .B2(new_n799), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n716), .A2(new_n442), .A3(new_n718), .A4(new_n777), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n789), .A2(new_n790), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n562), .A2(new_n426), .A3(G106gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n769), .A2(new_n770), .A3(new_n804), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n806), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n805), .A2(new_n806), .B1(new_n808), .B2(new_n802), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n542), .A2(new_n558), .A3(new_n548), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n549), .ZN(new_n813));
  INV_X1    g612(.A(new_n554), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n559), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n542), .A2(new_n548), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n550), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n811), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT55), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n813), .A2(new_n819), .A3(new_n822), .A4(new_n816), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n555), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n656), .B1(new_n655), .B2(new_n647), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n631), .A2(new_n632), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n634), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n644), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n660), .B2(new_n666), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n829), .A3(new_n685), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n824), .A2(new_n829), .A3(KEYINPUT114), .A4(new_n685), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n671), .A2(new_n824), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n829), .A2(new_n561), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n685), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n598), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n709), .A2(new_n672), .A3(new_n741), .A4(new_n562), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n689), .A3(new_n441), .A4(new_n443), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n672), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(G113gat), .Z(G1340gat));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n841), .A2(new_n562), .B1(new_n844), .B2(G120gat), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT116), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(KEYINPUT116), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n844), .A2(new_n846), .A3(G120gat), .A4(new_n847), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n846), .A2(new_n847), .B1(new_n844), .B2(G120gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  NOR2_X1   g649(.A1(new_n841), .A2(new_n598), .ZN(new_n851));
  XOR2_X1   g650(.A(KEYINPUT117), .B(G127gat), .Z(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1342gat));
  NOR2_X1   g652(.A1(new_n841), .A2(new_n741), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n855));
  AND2_X1   g654(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n854), .B2(new_n855), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(new_n598), .C1(new_n834), .C2(new_n837), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n839), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n442), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n840), .A2(new_n859), .A3(new_n442), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n702), .A2(new_n369), .A3(new_n692), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n867), .A3(new_n672), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT120), .B1(new_n868), .B2(new_n318), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n840), .A2(new_n870), .A3(new_n689), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n702), .A2(new_n426), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n840), .A2(new_n689), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n692), .B1(new_n874), .B2(KEYINPUT119), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n873), .A2(new_n318), .A3(new_n875), .A4(new_n671), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n868), .B2(new_n318), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n869), .A2(new_n877), .A3(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI221_X1 g678(.A(new_n876), .B1(KEYINPUT120), .B2(new_n879), .C1(new_n868), .C2(new_n318), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n315), .A3(new_n875), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n562), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(KEYINPUT121), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n882), .A2(new_n885), .A3(new_n562), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n864), .A2(new_n867), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n315), .C1(new_n887), .C2(new_n561), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n838), .A2(new_n839), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n426), .ZN(new_n891));
  INV_X1    g690(.A(new_n839), .ZN(new_n892));
  INV_X1    g691(.A(new_n837), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n709), .B1(new_n893), .B2(new_n830), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n859), .B(new_n442), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n891), .A2(new_n561), .A3(new_n866), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n889), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n884), .A2(new_n886), .B1(new_n888), .B2(new_n897), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n873), .A2(new_n875), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT123), .B1(new_n899), .B2(new_n598), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n873), .A2(new_n901), .A3(new_n875), .A4(new_n709), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n321), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n887), .A2(G155gat), .A3(new_n709), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  OAI21_X1  g704(.A(new_n322), .B1(new_n899), .B2(new_n741), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n741), .A2(new_n322), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n441), .A2(new_n689), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n840), .A2(new_n443), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n672), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n890), .B2(new_n689), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n840), .A2(KEYINPUT124), .A3(new_n369), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n914), .A2(new_n692), .A3(new_n443), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n671), .A2(new_n236), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n911), .A2(new_n237), .A3(new_n562), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n916), .A2(new_n562), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n237), .ZN(G1349gat));
  OAI21_X1  g720(.A(new_n229), .B1(new_n911), .B2(new_n598), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n709), .B1(new_n205), .B2(new_n204), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g724(.A1(new_n911), .A2(new_n741), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(G190gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n926), .B2(G190gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n685), .A2(new_n217), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n916), .B2(new_n930), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n891), .A2(new_n895), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n701), .A2(new_n910), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT125), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n672), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n914), .A2(new_n692), .A3(new_n872), .A4(new_n915), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n672), .A2(G197gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(new_n938), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n561), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n943), .A3(new_n561), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n938), .A2(G204gat), .A3(new_n562), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(new_n942), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n561), .A3(new_n935), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n945), .A2(new_n947), .A3(new_n950), .A4(new_n952), .ZN(G1353gat));
  OR3_X1    g752(.A1(new_n938), .A2(G211gat), .A3(new_n598), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n932), .A2(new_n709), .A3(new_n935), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n936), .A2(new_n959), .A3(new_n741), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n938), .B2(new_n741), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n963), .B(new_n959), .C1(new_n938), .C2(new_n741), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(G1355gat));
endmodule


