//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n204), .A2(G155gat), .A3(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT71), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n203), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT73), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT73), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n217), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT72), .B(new_n203), .C1(new_n205), .C2(new_n208), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n211), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n203), .ZN(new_n226));
  OAI22_X1  g025(.A1(new_n213), .A2(new_n215), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  AND2_X1   g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(KEYINPUT22), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G211gat), .B(G218gat), .Z(new_n233));
  XOR2_X1   g032(.A(new_n232), .B(new_n233), .Z(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n238), .A3(new_n227), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT68), .B(KEYINPUT29), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n235), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n235), .B2(new_n242), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(new_n229), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n244), .A2(new_n245), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G78gat), .B(G106gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G22gat), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT31), .B(G50gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n248), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254));
  XNOR2_X1  g053(.A(G8gat), .B(G36gat), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT70), .B(G64gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  AND2_X1   g061(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT27), .B(G183gat), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT65), .A3(KEYINPUT28), .A4(new_n262), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT26), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n276), .A2(new_n277), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n273), .A3(new_n274), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n262), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT24), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n295), .A3(new_n291), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n261), .B1(new_n297), .B2(new_n236), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n290), .A2(new_n295), .A3(new_n291), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n290), .B2(new_n291), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n260), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n235), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n261), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n241), .B1(new_n301), .B2(new_n279), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n234), .B(new_n304), .C1(new_n305), .C2(new_n261), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT69), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT69), .B1(new_n303), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n259), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(new_n259), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(KEYINPUT30), .A3(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n312), .A2(KEYINPUT30), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT66), .B1(new_n320), .B2(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(G113gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT67), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325));
  XOR2_X1   g124(.A(G127gat), .B(G134gat), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n328), .B(new_n319), .C1(new_n321), .C2(new_n322), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n318), .A2(G120gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n325), .B1(new_n331), .B2(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n224), .A2(new_n330), .A3(new_n333), .A4(new_n227), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n329), .A2(new_n325), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n326), .B1(new_n323), .B2(KEYINPUT67), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(new_n332), .B2(new_n326), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n227), .A4(new_n224), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n330), .A2(new_n333), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n240), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n342), .A2(KEYINPUT74), .A3(new_n343), .A4(new_n240), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n316), .B(new_n341), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n334), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n227), .A2(new_n224), .B1(new_n330), .B2(new_n333), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n316), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n228), .A2(new_n343), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n315), .B1(new_n354), .B2(new_n334), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(new_n358), .A3(KEYINPUT5), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n346), .A2(new_n347), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(new_n315), .A3(new_n336), .A4(new_n340), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT77), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n364), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n359), .A2(new_n364), .A3(new_n374), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n372), .ZN(new_n378));
  AOI221_X4 g177(.A(new_n254), .B1(new_n313), .B2(new_n314), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n378), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n313), .A2(new_n314), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT78), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n253), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G15gat), .B(G43gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(G227gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n297), .A2(new_n343), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n301), .A2(new_n339), .A3(new_n279), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n386), .B1(new_n391), .B2(KEYINPUT33), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT34), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n390), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(G227gat), .A3(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n389), .B(new_n390), .C1(new_n387), .C2(new_n388), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n394), .B2(new_n398), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n392), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n398), .ZN(new_n404));
  INV_X1    g203(.A(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n392), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n400), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT36), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n412), .A2(KEYINPUT39), .A3(new_n315), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n374), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n354), .A2(new_n315), .A3(new_n334), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT39), .B(new_n415), .C1(new_n412), .C2(new_n315), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n414), .A2(KEYINPUT40), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT40), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n417), .A2(new_n418), .A3(new_n377), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n381), .A2(KEYINPUT79), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n313), .A2(new_n421), .A3(new_n314), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n253), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT37), .B1(new_n303), .B2(new_n306), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(new_n259), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n298), .A2(new_n302), .A3(new_n235), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n304), .B1(new_n305), .B2(new_n261), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n235), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT37), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n425), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n311), .B1(new_n438), .B2(new_n428), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT81), .A3(new_n426), .A4(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n312), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n375), .A2(KEYINPUT82), .A3(new_n371), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n259), .B1(new_n429), .B2(new_n430), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n307), .A2(new_n308), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT38), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n370), .A2(new_n371), .A3(new_n375), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT82), .B1(new_n375), .B2(new_n371), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n443), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n423), .B(new_n424), .C1(new_n442), .C2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n383), .A2(new_n411), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n374), .B1(new_n359), .B2(new_n364), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n377), .A2(new_n454), .A3(new_n372), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n375), .A2(new_n373), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n381), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n254), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n409), .A2(new_n253), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n409), .B1(new_n420), .B2(new_n422), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n461), .A2(KEYINPUT35), .B1(new_n465), .B2(new_n424), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n453), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n468));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n469));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NOR3_X1   g273(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(G29gat), .A2(G36gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n469), .B2(new_n470), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n475), .B(KEYINPUT85), .Z(new_n482));
  OAI221_X1 g281(.A(new_n481), .B1(new_n470), .B2(new_n469), .C1(new_n482), .C2(new_n474), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  OAI221_X1 g287(.A(new_n487), .B1(KEYINPUT86), .B2(new_n488), .C1(G1gat), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n489), .B(new_n490), .Z(new_n491));
  OR3_X1    g290(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT87), .B1(new_n484), .B2(new_n491), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n480), .A2(new_n483), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n468), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n494), .A2(new_n497), .A3(KEYINPUT18), .A4(new_n499), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n492), .A2(KEYINPUT88), .A3(new_n493), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n504), .A2(new_n505), .B1(new_n484), .B2(new_n491), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n499), .B(KEYINPUT13), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n501), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  INV_X1    g308(.A(G197gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT11), .B(G169gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT12), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n484), .A2(new_n491), .ZN(new_n517));
  INV_X1    g316(.A(new_n505), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT88), .B1(new_n492), .B2(new_n493), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n507), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(new_n514), .A3(new_n501), .A4(new_n502), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n202), .B1(new_n467), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT89), .B(new_n524), .C1(new_n453), .C2(new_n466), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g333(.A(G99gat), .ZN(new_n535));
  INV_X1    g334(.A(G106gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT8), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n534), .B(new_n537), .C1(G85gat), .C2(G92gat), .ZN(new_n538));
  XOR2_X1   g337(.A(G99gat), .B(G106gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n532), .B1(new_n484), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n496), .A2(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n531), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n531), .A2(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  OR2_X1    g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n562));
  INV_X1    g361(.A(new_n559), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n491), .B1(new_n556), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT91), .Z(new_n569));
  INV_X1    g368(.A(G127gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n556), .ZN(new_n572));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n569), .B(G127gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G155gat), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n577), .B2(new_n580), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n540), .B(new_n567), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT95), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n540), .A2(new_n567), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT10), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g399(.A(KEYINPUT94), .B(new_n592), .C1(new_n595), .C2(new_n597), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n589), .B(new_n594), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n588), .B1(new_n598), .B2(new_n593), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n555), .A2(new_n585), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n528), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n380), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g412(.A1(new_n420), .A2(new_n422), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT16), .B(G8gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT42), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT98), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  AOI211_X1 g418(.A(new_n614), .B(new_n619), .C1(new_n608), .C2(new_n609), .ZN(new_n620));
  INV_X1    g419(.A(new_n614), .ZN(new_n621));
  AOI21_X1  g420(.A(G8gat), .B1(new_n610), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n622), .B2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g422(.A(new_n409), .ZN(new_n624));
  AOI21_X1  g423(.A(G15gat), .B1(new_n610), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n411), .B1(new_n608), .B2(new_n609), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(G15gat), .B2(new_n626), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n253), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  INV_X1    g429(.A(new_n555), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n585), .A2(new_n604), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n528), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n633), .A2(G29gat), .A3(new_n380), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT45), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n516), .A2(new_n523), .A3(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT99), .B1(new_n516), .B2(new_n523), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n632), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n465), .A2(new_n424), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n383), .A2(new_n411), .A3(new_n452), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n555), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT100), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n631), .B1(new_n453), .B2(new_n466), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT44), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n555), .A2(KEYINPUT44), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n453), .A2(new_n466), .A3(KEYINPUT101), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n645), .B2(new_n646), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n654), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n642), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G29gat), .B1(new_n660), .B2(new_n380), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n635), .A2(new_n661), .ZN(G1328gat));
  NOR3_X1   g461(.A1(new_n633), .A2(G36gat), .A3(new_n614), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT46), .ZN(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n660), .B2(new_n614), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(G43gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n411), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n633), .A2(G43gat), .A3(new_n409), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT47), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n648), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n651), .B1(new_n650), .B2(KEYINPUT44), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n658), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n668), .A3(new_n641), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(KEYINPUT102), .A3(G43gat), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(KEYINPUT47), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n555), .B(new_n640), .C1(new_n526), .C2(new_n527), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n667), .A3(new_n624), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n680), .A2(new_n683), .A3(new_n667), .A4(new_n624), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n671), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT104), .B(new_n671), .C1(new_n679), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1330gat));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  INV_X1    g490(.A(G50gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n680), .A2(new_n692), .A3(new_n253), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT105), .Z(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n659), .B2(new_n253), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n698), .B(KEYINPUT48), .C1(new_n697), .C2(new_n693), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(G1331gat));
  NOR2_X1   g499(.A1(new_n655), .A2(new_n657), .ZN(new_n701));
  INV_X1    g500(.A(new_n585), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n631), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n524), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n636), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n605), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n380), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT107), .B(G57gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  NOR2_X1   g512(.A1(new_n710), .A2(new_n614), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  AND2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n715), .ZN(G1333gat));
  AND2_X1   g517(.A1(new_n705), .A2(new_n709), .ZN(new_n719));
  INV_X1    g518(.A(G71gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n624), .ZN(new_n721));
  OAI21_X1  g520(.A(G71gat), .B1(new_n710), .B2(new_n411), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT108), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n724), .A2(KEYINPUT50), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n719), .A2(new_n253), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n708), .A2(new_n585), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n647), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n737), .B(new_n738), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n604), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n611), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n605), .B1(new_n653), .B2(new_n658), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n734), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n743), .A3(new_n734), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n380), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n742), .B1(new_n748), .B2(G85gat), .ZN(G1336gat));
  NOR3_X1   g548(.A1(new_n740), .A2(G92gat), .A3(new_n614), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n744), .A2(new_n734), .ZN(new_n753));
  OAI21_X1  g552(.A(G92gat), .B1(new_n753), .B2(new_n614), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n747), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n621), .B1(new_n756), .B2(new_n745), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n750), .B1(new_n757), .B2(G92gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n752), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n535), .A3(new_n624), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n411), .B1(new_n746), .B2(new_n747), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n535), .ZN(G1338gat));
  NOR3_X1   g561(.A1(new_n740), .A2(G106gat), .A3(new_n424), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G106gat), .B1(new_n753), .B2(new_n424), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n253), .B1(new_n756), .B2(new_n745), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n763), .B1(new_n768), .B2(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n606), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n772), .B2(new_n708), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n639), .A2(new_n606), .A3(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n595), .A2(new_n597), .A3(new_n592), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n778), .B(KEYINPUT54), .C1(new_n600), .C2(new_n601), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n780));
  NAND2_X1  g579(.A1(new_n598), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n588), .A4(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n602), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n588), .A3(new_n781), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n786), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n506), .A2(new_n507), .B1(new_n500), .B2(new_n498), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(new_n513), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n523), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n631), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(new_n605), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n793), .B2(new_n708), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n777), .B(new_n798), .C1(new_n800), .C2(new_n631), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n702), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n784), .A2(new_n602), .A3(new_n785), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n790), .A2(new_n792), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n803), .B(new_n804), .C1(new_n637), .C2(new_n638), .ZN(new_n805));
  INV_X1    g604(.A(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n555), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n777), .B1(new_n808), .B2(new_n798), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n776), .B1(new_n802), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n380), .A2(new_n253), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n462), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n525), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n708), .A2(new_n318), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(G1340gat));
  NAND4_X1  g614(.A1(new_n810), .A2(new_n462), .A3(new_n604), .A4(new_n811), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n320), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n822));
  NOR4_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n818), .A4(new_n320), .ZN(new_n823));
  INV_X1    g622(.A(new_n822), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(new_n820), .B1(KEYINPUT117), .B2(G120gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n823), .A2(new_n825), .ZN(G1341gat));
  AND2_X1   g625(.A1(KEYINPUT119), .A2(G127gat), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT119), .A2(G127gat), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n702), .ZN(new_n830));
  MUX2_X1   g629(.A(new_n827), .B(new_n829), .S(new_n830), .Z(G1342gat));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n462), .A3(new_n631), .A4(new_n811), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G134gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(G134gat), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n835), .A2(KEYINPUT120), .A3(new_n834), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT120), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  OAI221_X1 g636(.A(new_n833), .B1(new_n834), .B2(new_n835), .C1(new_n836), .C2(new_n837), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n668), .A2(new_n380), .A3(new_n621), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n810), .B2(new_n253), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n524), .A2(new_n789), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n786), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n555), .B1(new_n844), .B2(new_n799), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n585), .B1(new_n845), .B2(new_n798), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n776), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n253), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n773), .A2(new_n775), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n253), .C1(new_n850), .C2(new_n846), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n840), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n212), .B1(new_n855), .B2(new_n524), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n810), .A2(new_n253), .ZN(new_n857));
  NOR4_X1   g656(.A1(new_n857), .A2(G141gat), .A3(new_n525), .A4(new_n840), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT58), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n849), .A2(new_n853), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n708), .B(new_n839), .C1(new_n841), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n858), .B1(new_n861), .B2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n856), .A2(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n857), .A2(new_n840), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n214), .A3(new_n604), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n604), .B(new_n839), .C1(new_n841), .C2(new_n860), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(G148gat), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n606), .A2(new_n525), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n871), .B(new_n253), .C1(new_n846), .C2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n870), .A2(new_n604), .A3(new_n839), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n868), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n866), .B1(new_n869), .B2(new_n876), .ZN(G1345gat));
  AOI21_X1  g676(.A(G155gat), .B1(new_n865), .B2(new_n585), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n702), .A2(new_n206), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n855), .B2(new_n879), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n865), .B2(new_n631), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n555), .A2(new_n207), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n855), .B2(new_n882), .ZN(G1347gat));
  INV_X1    g682(.A(new_n460), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n631), .B1(new_n805), .B2(new_n806), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n793), .A2(new_n631), .A3(new_n797), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT116), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n702), .A3(new_n801), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(new_n776), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n611), .A2(new_n614), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n525), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n708), .A2(new_n273), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(G1348gat));
  NOR2_X1   g693(.A1(new_n891), .A2(new_n605), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(new_n274), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n889), .A2(new_n585), .A3(new_n890), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n270), .B1(new_n898), .B2(G183gat), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n897), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n898), .A2(new_n284), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT60), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n900), .B(new_n906), .C1(new_n901), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1350gat));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G190gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n555), .ZN(new_n911));
  MUX2_X1   g710(.A(new_n909), .B(new_n910), .S(new_n911), .Z(G1351gat));
  INV_X1    g711(.A(new_n874), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n857), .B2(KEYINPUT57), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n890), .A2(new_n411), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n914), .A2(new_n915), .A3(new_n524), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n424), .B1(new_n888), .B2(new_n776), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n874), .B(new_n917), .C1(new_n919), .C2(new_n871), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT125), .B1(new_n920), .B2(new_n525), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n921), .A3(G197gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n810), .A2(new_n253), .A3(new_n917), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(KEYINPUT123), .A3(new_n917), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n510), .A3(new_n708), .A4(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n932), .A3(new_n917), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n933), .A2(new_n605), .B1(new_n934), .B2(KEYINPUT62), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(KEYINPUT126), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n934), .B(KEYINPUT62), .C1(new_n933), .C2(new_n605), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n914), .A2(new_n604), .A3(new_n917), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n932), .C2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n914), .A2(new_n585), .A3(new_n917), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n942));
  OAI211_X1 g741(.A(KEYINPUT63), .B(G211gat), .C1(new_n920), .C2(new_n702), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n926), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n702), .A2(G211gat), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n942), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  NAND4_X1  g746(.A1(new_n870), .A2(KEYINPUT127), .A3(new_n874), .A4(new_n917), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n920), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n948), .A2(new_n950), .A3(new_n631), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G218gat), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n945), .A2(G218gat), .A3(new_n555), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1355gat));
endmodule


