//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT69), .B(G113gat), .Z(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n202), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n208), .B(KEYINPUT67), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n202), .A2(G113gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(KEYINPUT1), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT71), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n219), .A2(KEYINPUT24), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .B1(new_n220), .B2(KEYINPUT24), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT25), .B1(new_n224), .B2(KEYINPUT64), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n223), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n225), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n222), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n227), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(new_n220), .C1(new_n232), .C2(new_n231), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT28), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n238), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n230), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n218), .B(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G15gat), .B(G43gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT33), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(KEYINPUT32), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT73), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(KEYINPUT32), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n247), .A2(new_n257), .A3(KEYINPUT32), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n250), .B1(new_n247), .B2(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n245), .A2(new_n246), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT34), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n254), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n262), .B(KEYINPUT34), .Z(new_n265));
  OR2_X1    g064(.A1(new_n253), .A2(KEYINPUT73), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n253), .A2(KEYINPUT73), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n264), .A2(new_n269), .A3(KEYINPUT36), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n256), .A2(new_n259), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT74), .B1(new_n272), .B2(new_n265), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n274), .B(new_n263), .C1(new_n254), .C2(new_n261), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n265), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n277), .B2(KEYINPUT36), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279));
  INV_X1    g078(.A(G155gat), .ZN(new_n280));
  INV_X1    g079(.A(G162gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT2), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT79), .ZN(new_n283));
  XNOR2_X1  g082(.A(G155gat), .B(G162gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n284), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n284), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(KEYINPUT2), .B2(new_n285), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n215), .A3(new_n211), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n218), .A2(new_n293), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n293), .A2(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n216), .ZN(new_n304));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n296), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n306), .B(new_n308), .C1(new_n298), .C2(new_n296), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n216), .A2(new_n293), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n305), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT81), .ZN(new_n316));
  XOR2_X1   g115(.A(G57gat), .B(G85gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n307), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n307), .A2(new_n314), .A3(KEYINPUT82), .A4(new_n321), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(new_n307), .B2(new_n314), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT6), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340));
  OAI22_X1  g139(.A1(new_n338), .A2(KEYINPUT22), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(KEYINPUT75), .ZN(new_n343));
  NOR2_X1   g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n343), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n244), .B(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AND4_X1   g150(.A1(G226gat), .A2(new_n230), .A3(G233gat), .A4(new_n243), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(G226gat), .A3(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n346), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n244), .A2(new_n349), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n353), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n354), .B1(new_n353), .B2(new_n358), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n336), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n358), .A3(new_n335), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n279), .B1(new_n332), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n346), .B1(new_n302), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n346), .A2(new_n368), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n294), .B1(new_n370), .B2(new_n301), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n345), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n374), .B2(new_n341), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n342), .A2(new_n345), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT3), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n294), .B2(new_n377), .ZN(new_n378));
  OAI22_X1  g177(.A1(new_n372), .A2(new_n373), .B1(new_n369), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT31), .B(G50gat), .Z(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G22gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n381), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n365), .A2(new_n364), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n329), .A2(new_n331), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT83), .A4(new_n361), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n353), .A2(new_n358), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT37), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n391), .A2(KEYINPUT38), .A3(new_n335), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  OAI221_X1 g192(.A(new_n356), .B1(new_n244), .B2(new_n393), .C1(new_n348), .C2(new_n350), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n355), .A2(new_n357), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT85), .B(new_n394), .C1(new_n395), .C2(new_n356), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT37), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n351), .A2(new_n346), .A3(new_n352), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n396), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n329), .A2(new_n331), .A3(new_n362), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n360), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n353), .A2(new_n358), .A3(new_n354), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n398), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT87), .B1(new_n409), .B2(new_n335), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT37), .B1(new_n359), .B2(new_n360), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n336), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n410), .B(new_n413), .C1(KEYINPUT37), .C2(new_n390), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n414), .B2(KEYINPUT38), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n305), .B1(new_n299), .B2(new_n304), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT39), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT39), .B1(new_n311), .B2(new_n312), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n418), .B(new_n321), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n330), .B1(new_n421), .B2(KEYINPUT40), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n366), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT40), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n420), .A2(KEYINPUT84), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT84), .B1(new_n420), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n384), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n278), .B(new_n389), .C1(new_n415), .C2(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n332), .A2(new_n366), .A3(KEYINPUT35), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n264), .A2(new_n385), .A3(new_n269), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n273), .A2(new_n384), .A3(new_n275), .A4(new_n276), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n367), .B2(new_n388), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT35), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT16), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(G1gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(G1gat), .B2(new_n438), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G8gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G29gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT14), .B(G29gat), .Z(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(G36gat), .ZN(new_n447));
  XOR2_X1   g246(.A(G43gat), .B(G50gat), .Z(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT88), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n450));
  XNOR2_X1  g249(.A(G43gat), .B(G50gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(new_n450), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n447), .A2(new_n455), .B1(new_n449), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT17), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n447), .A2(new_n455), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n449), .A2(new_n453), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n443), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n454), .A2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n463), .A2(KEYINPUT18), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n464), .B(KEYINPUT13), .Z(new_n468));
  INV_X1    g267(.A(new_n466), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n442), .A2(new_n465), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G197gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT11), .B(G169gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT12), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n467), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT18), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n471), .A3(new_n467), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n437), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G71gat), .A2(G78gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(G71gat), .A2(G78gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494));
  NAND3_X1  g293(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT92), .ZN(new_n500));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n496), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G57gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(KEYINPUT93), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(G57gat), .ZN(new_n507));
  OAI21_X1  g306(.A(G64gat), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n499), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G64gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n490), .A2(new_n493), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G183gat), .B(G211gat), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n517), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n516), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n514), .A2(KEYINPUT96), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n502), .A2(new_n527), .A3(new_n513), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(KEYINPUT21), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n529), .A2(new_n443), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n529), .B2(new_n443), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n525), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n520), .A3(new_n524), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G190gat), .B(G218gat), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(G99gat), .B2(G106gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT8), .ZN(new_n552));
  OR2_X1    g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT97), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n545), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G99gat), .B(G106gat), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT99), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT7), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n553), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT97), .B1(new_n552), .B2(new_n553), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n557), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT98), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n554), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n557), .A4(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n565), .A2(new_n566), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n566), .B1(new_n565), .B2(new_n572), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n542), .B1(new_n575), .B2(new_n465), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n565), .A2(new_n572), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT100), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n558), .A2(new_n564), .B1(new_n568), .B2(new_n571), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n566), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n457), .A2(new_n462), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n577), .B(new_n583), .C1(new_n573), .C2(new_n574), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n541), .B(new_n576), .C1(new_n584), .C2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n583), .B1(new_n573), .B2(new_n574), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT101), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n585), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n541), .B1(new_n591), .B2(new_n576), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n588), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n576), .B1(new_n584), .B2(new_n586), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n540), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n599), .B2(new_n587), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n539), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n596), .B1(new_n588), .B2(new_n592), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n595), .A3(new_n587), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n539), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT103), .ZN(new_n610));
  INV_X1    g409(.A(new_n528), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n527), .B1(new_n502), .B2(new_n513), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n579), .A2(new_n581), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n514), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n562), .A2(new_n556), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n572), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n618), .B(new_n613), .C1(new_n616), .C2(new_n580), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n610), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n610), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n578), .A2(new_n514), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(new_n618), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n620), .A2(new_n623), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n489), .A2(new_n608), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n332), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g434(.A1(new_n608), .A2(new_n632), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n437), .A2(new_n366), .A3(new_n488), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT42), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT105), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n637), .A2(KEYINPUT104), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(KEYINPUT104), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(G8gat), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n638), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n641), .B(new_n644), .C1(KEYINPUT42), .C2(new_n646), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n264), .A2(new_n269), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n278), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n652), .B2(new_n648), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n489), .A2(new_n384), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n636), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT106), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n657), .A3(new_n636), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n656), .B2(new_n658), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n606), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n278), .A2(new_n389), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n413), .B1(KEYINPUT37), .B2(new_n390), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n412), .B1(new_n411), .B2(new_n336), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT38), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n406), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n428), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n433), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n367), .A2(new_n388), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n673), .A2(KEYINPUT35), .B1(new_n431), .B2(new_n430), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n663), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n437), .A2(KEYINPUT44), .A3(new_n663), .ZN(new_n678));
  INV_X1    g477(.A(new_n488), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n632), .A2(new_n679), .A3(new_n539), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n677), .A2(new_n332), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G29gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n632), .A2(new_n539), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n663), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n387), .A2(G29gat), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n437), .A2(new_n488), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n682), .A2(new_n689), .A3(KEYINPUT108), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1328gat));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n366), .A3(new_n678), .A4(new_n680), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G36gat), .ZN(new_n696));
  INV_X1    g495(.A(new_n366), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(G36gat), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n437), .A2(new_n488), .A3(new_n685), .A4(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(new_n701), .A3(KEYINPUT109), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n677), .A2(new_n651), .A3(new_n678), .A4(new_n680), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n649), .ZN(new_n709));
  OR4_X1    g508(.A1(G43gat), .A2(new_n489), .A3(new_n709), .A4(new_n684), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n708), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1330gat));
  NAND4_X1  g513(.A1(new_n677), .A2(new_n385), .A3(new_n678), .A4(new_n680), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n654), .A2(new_n717), .A3(new_n685), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  NOR3_X1   g522(.A1(new_n608), .A2(new_n488), .A3(new_n631), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n437), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n387), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT93), .B(G57gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT49), .B(G64gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n366), .A3(new_n730), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n725), .A2(new_n697), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT110), .Z(G1333gat));
  NOR3_X1   g533(.A1(new_n725), .A2(G71gat), .A3(new_n709), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n651), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(G71gat), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n729), .A2(new_n385), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n631), .A2(new_n488), .A3(new_n539), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n677), .A2(new_n678), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n387), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n606), .B1(new_n429), .B2(new_n436), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n488), .A2(new_n539), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n744), .A2(KEYINPUT51), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n387), .A2(G85gat), .A3(new_n631), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT111), .Z(new_n750));
  OAI21_X1  g549(.A(new_n743), .B1(new_n748), .B2(new_n750), .ZN(G1336gat));
  NAND4_X1  g550(.A1(new_n677), .A2(new_n366), .A3(new_n678), .A4(new_n741), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n697), .A2(G92gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n632), .B(new_n754), .C1(new_n746), .C2(new_n747), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n742), .B2(new_n278), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n709), .A2(G99gat), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n632), .B(new_n762), .C1(new_n746), .C2(new_n747), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1338gat));
  NAND4_X1  g563(.A1(new_n677), .A2(new_n385), .A3(new_n678), .A4(new_n741), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n384), .A2(G106gat), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n632), .B(new_n767), .C1(new_n746), .C2(new_n747), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n766), .A2(new_n768), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1339gat));
  NAND4_X1  g573(.A1(new_n603), .A2(new_n679), .A3(new_n607), .A4(new_n631), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n469), .A2(new_n470), .A3(new_n468), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n475), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n484), .B(new_n779), .C1(new_n628), .C2(new_n630), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT113), .Z(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n615), .A2(new_n619), .A3(new_n610), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n783), .A2(new_n620), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n619), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n526), .A2(KEYINPUT10), .A3(new_n528), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n573), .A2(new_n574), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(new_n621), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n629), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n782), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n630), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n621), .B1(new_n786), .B2(new_n788), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n615), .A2(new_n619), .A3(new_n610), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n627), .B1(new_n620), .B2(new_n784), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n791), .A2(new_n488), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n606), .B1(new_n781), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n791), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n792), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n484), .A2(new_n779), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n606), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n539), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n776), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n385), .A3(new_n709), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n366), .A2(new_n387), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n679), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n808), .A2(new_n387), .A3(new_n433), .A4(new_n366), .ZN(new_n813));
  INV_X1    g612(.A(new_n206), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n488), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1340gat));
  NOR3_X1   g615(.A1(new_n811), .A2(new_n202), .A3(new_n631), .ZN(new_n817));
  AOI21_X1  g616(.A(G120gat), .B1(new_n813), .B2(new_n632), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  OAI21_X1  g618(.A(G127gat), .B1(new_n811), .B2(new_n807), .ZN(new_n820));
  INV_X1    g619(.A(G127gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n821), .A3(new_n539), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1342gat));
  INV_X1    g622(.A(G134gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n813), .A2(new_n824), .A3(new_n663), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n811), .B2(new_n606), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n808), .B2(new_n384), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT115), .B(new_n831), .C1(new_n808), .C2(new_n384), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n384), .A2(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n798), .A2(new_n780), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n663), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n798), .A2(KEYINPUT116), .A3(new_n780), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n807), .B1(new_n841), .B2(new_n804), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n836), .B1(new_n843), .B2(new_n776), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n834), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n278), .A2(new_n810), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n488), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n278), .A2(new_n385), .ZN(new_n850));
  NOR4_X1   g649(.A1(new_n850), .A2(new_n808), .A3(new_n387), .A4(new_n366), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n288), .A3(new_n488), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(G148gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n851), .A2(new_n858), .A3(new_n632), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n846), .A2(new_n632), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n806), .A2(new_n807), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n775), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n836), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT102), .B1(new_n606), .B2(new_n539), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n602), .B(new_n807), .C1(new_n604), .C2(new_n605), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n679), .A4(new_n631), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n775), .A2(KEYINPUT117), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n804), .B1(new_n839), .B2(new_n840), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n539), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n384), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n870), .A4(new_n869), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n876), .B2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n878), .B(KEYINPUT57), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n861), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n860), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n845), .A2(new_n632), .A3(new_n846), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n858), .A2(KEYINPUT59), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n859), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT120), .B(new_n859), .C1(new_n881), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n851), .A2(new_n280), .A3(new_n539), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n847), .A2(new_n539), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n280), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n851), .B2(new_n663), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n606), .A2(new_n281), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n847), .B2(new_n894), .ZN(G1347gat));
  INV_X1    g694(.A(G169gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n697), .A2(new_n332), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n809), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n488), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT122), .Z(new_n900));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n387), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT121), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n433), .A2(new_n697), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n896), .A3(new_n488), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(G1348gat));
  INV_X1    g705(.A(G176gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n907), .A3(new_n632), .ZN(new_n908));
  INV_X1    g707(.A(new_n898), .ZN(new_n909));
  OAI21_X1  g708(.A(G176gat), .B1(new_n909), .B2(new_n631), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1349gat));
  NOR2_X1   g710(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n902), .A2(new_n236), .A3(new_n539), .A4(new_n903), .ZN(new_n913));
  OAI21_X1  g712(.A(G183gat), .B1(new_n909), .B2(new_n807), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n915), .B(new_n916), .Z(G1350gat));
  AOI21_X1  g716(.A(new_n237), .B1(new_n898), .B2(new_n663), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT61), .Z(new_n919));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n237), .A3(new_n663), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n850), .A2(new_n697), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n902), .ZN(new_n924));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n488), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n278), .A2(new_n897), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n874), .A2(new_n875), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n878), .B1(new_n927), .B2(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n864), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT125), .B1(new_n877), .B2(new_n879), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n488), .A2(G197gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n631), .A2(G204gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n923), .A2(new_n902), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT62), .Z(new_n938));
  NAND3_X1  g737(.A1(new_n278), .A2(new_n632), .A3(new_n897), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n931), .B2(new_n932), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n923), .A2(new_n945), .A3(new_n539), .A4(new_n902), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n877), .A2(new_n879), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n278), .A2(new_n539), .A3(new_n897), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n951), .A2(KEYINPUT63), .A3(new_n945), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(new_n945), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n952), .A3(new_n953), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n924), .B2(new_n663), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n663), .A2(G218gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n933), .B2(new_n956), .ZN(G1355gat));
endmodule


