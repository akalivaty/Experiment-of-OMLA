//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT75), .B(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT76), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(KEYINPUT76), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  XOR2_X1   g020(.A(G155gat), .B(G162gat), .Z(new_n222));
  AOI22_X1  g021(.A1(new_n211), .A2(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(G211gat), .ZN(new_n227));
  INV_X1    g026(.A(G218gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(KEYINPUT22), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n224), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n217), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n222), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n236), .A2(new_n237), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n232), .B(KEYINPUT72), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n245), .B2(new_n225), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G228gat), .A3(G233gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT31), .B(G50gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n244), .B2(new_n247), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n204), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n203), .A3(new_n250), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT27), .B(G183gat), .Z(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G190gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(G190gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n259), .A2(KEYINPUT67), .B1(new_n260), .B2(KEYINPUT28), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(KEYINPUT67), .B2(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G169gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n267), .A2(KEYINPUT26), .A3(new_n268), .ZN(new_n269));
  AOI211_X1 g068(.A(new_n264), .B(new_n269), .C1(KEYINPUT26), .C2(new_n268), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(KEYINPUT23), .B2(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(KEYINPUT23), .B2(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n278), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n280), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n288), .A3(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(new_n245), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  AND2_X1   g096(.A1(new_n285), .A2(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n290), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n294), .B(new_n297), .C1(new_n300), .C2(new_n232), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT73), .B1(new_n271), .B2(new_n284), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n288), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n289), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n233), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n310), .A2(KEYINPUT74), .A3(new_n294), .A4(new_n297), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n294), .A4(new_n297), .ZN(new_n313));
  INV_X1    g112(.A(new_n297), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n232), .B1(new_n307), .B2(new_n308), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  OR3_X1    g124(.A1(new_n323), .A2(new_n325), .A3(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT1), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n324), .A2(new_n326), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n327), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n322), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n223), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n331), .A2(new_n333), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n241), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n241), .A2(new_n336), .A3(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n223), .A2(new_n224), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n336), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n335), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n340), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G1gat), .B(G29gat), .Z(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n341), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n339), .A2(new_n342), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(KEYINPUT39), .C1(new_n341), .C2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n359), .C1(KEYINPUT39), .C2(new_n363), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT40), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n367), .B2(new_n366), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n312), .A2(new_n318), .A3(KEYINPUT82), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n321), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT37), .B1(new_n315), .B2(new_n316), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n314), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT37), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n294), .C1(new_n300), .C2(new_n232), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n310), .A2(KEYINPUT85), .A3(new_n376), .A4(new_n294), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n372), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT87), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n374), .B1(new_n379), .B2(new_n380), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n314), .A2(new_n372), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n291), .A2(new_n292), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n389), .A2(new_n293), .B1(new_n309), .B2(new_n233), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n390), .B2(KEYINPUT37), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n303), .A2(new_n311), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT80), .B1(new_n361), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n351), .A2(new_n353), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n351), .B2(new_n344), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n400));
  INV_X1    g199(.A(new_n396), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n360), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n352), .A2(new_n354), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n359), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n361), .A3(new_n396), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n405), .A2(KEYINPUT83), .A3(new_n361), .A4(new_n396), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n381), .A2(new_n391), .A3(KEYINPUT86), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n256), .B(new_n371), .C1(new_n387), .C2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G71gat), .B(G99gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT70), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(KEYINPUT70), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT33), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n285), .B(new_n334), .ZN(new_n420));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n421), .B(KEYINPUT64), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI221_X1 g222(.A(KEYINPUT32), .B1(new_n417), .B2(new_n419), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n420), .A2(new_n423), .B1(KEYINPUT32), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n426), .A2(new_n427), .A3(new_n416), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n426), .B2(new_n416), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(new_n431), .A3(new_n423), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n421), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT34), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n420), .A2(KEYINPUT71), .A3(new_n431), .A4(new_n423), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n438), .B(new_n424), .C1(new_n429), .C2(new_n428), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT36), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n253), .A2(new_n255), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n406), .A2(new_n402), .A3(new_n397), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n319), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n440), .A2(new_n256), .A3(new_n441), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n319), .A2(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n321), .A2(new_n370), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n410), .A2(KEYINPUT35), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n413), .A2(new_n451), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT96), .ZN(new_n461));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(G197gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT11), .B(G169gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(G43gat), .A2(G50gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(G43gat), .A2(G50gat), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT15), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(KEYINPUT90), .A2(G29gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(KEYINPUT90), .A2(G29gat), .ZN(new_n476));
  OAI21_X1  g275(.A(G36gat), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n482));
  INV_X1    g281(.A(G36gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G43gat), .ZN(new_n489));
  INV_X1    g288(.A(G50gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n477), .A3(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n488), .A2(new_n495), .A3(KEYINPUT92), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n472), .A2(new_n477), .A3(new_n494), .ZN(new_n498));
  NOR4_X1   g297(.A1(KEYINPUT91), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n486), .B1(new_n482), .B2(new_n483), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n478), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n481), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT16), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n507), .A2(G1gat), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT93), .B(new_n506), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n514), .A2(new_n510), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n481), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT92), .B1(new_n488), .B2(new_n495), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n497), .A3(new_n501), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n518), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n503), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(KEYINPUT18), .A3(new_n525), .A4(new_n527), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n503), .A2(new_n526), .A3(KEYINPUT94), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n522), .B2(new_n518), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n522), .A2(new_n518), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n525), .B(KEYINPUT13), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n530), .A2(new_n468), .A3(new_n531), .A4(new_n538), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n531), .A2(new_n538), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(KEYINPUT95), .A3(new_n468), .A4(new_n530), .ZN(new_n544));
  AOI221_X4 g343(.A(new_n461), .B1(new_n469), .B2(new_n539), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(new_n469), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT96), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT20), .Z(new_n552));
  AOI21_X1  g351(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT97), .ZN(new_n554));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G57gat), .B(G64gat), .Z(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(new_n565), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n552), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  INV_X1    g369(.A(new_n552), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n518), .B1(new_n562), .B2(new_n561), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n574), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n569), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n575), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT99), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n586), .A2(KEYINPUT41), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n593), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n593), .A3(new_n599), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n592), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  INV_X1    g403(.A(new_n592), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n604), .A2(new_n605), .A3(new_n600), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n591), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n604), .B2(new_n600), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n601), .A2(new_n592), .A3(new_n602), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT101), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n611), .A2(new_n503), .B1(KEYINPUT41), .B2(new_n586), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT102), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n607), .A2(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n505), .A3(new_n523), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n612), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n590), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n589), .A3(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n561), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n607), .A2(new_n610), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n595), .A2(new_n599), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT103), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n558), .A3(new_n560), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n603), .B2(new_n606), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n609), .A3(new_n608), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT10), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G230gat), .ZN(new_n634));
  INV_X1    g433(.A(G233gat), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n626), .A2(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n636), .B2(new_n638), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g444(.A1(new_n583), .A2(new_n621), .A3(new_n623), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n460), .A2(new_n550), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n447), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n508), .ZN(G1324gat));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n456), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n506), .B2(new_n650), .ZN(new_n653));
  MUX2_X1   g452(.A(new_n652), .B(new_n653), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g453(.A1(new_n443), .A2(new_n445), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n647), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n442), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n647), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n647), .A2(new_n256), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n583), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n645), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n621), .A2(new_n623), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n312), .A2(new_n318), .A3(KEYINPUT82), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT82), .B1(new_n312), .B2(new_n318), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n446), .B1(new_n669), .B2(new_n369), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n410), .A2(new_n411), .A3(new_n395), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n671), .A2(new_n394), .A3(new_n386), .A4(new_n383), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n450), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n440), .A2(new_n256), .A3(new_n441), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(new_n457), .B1(new_n454), .B2(KEYINPUT35), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n550), .B(new_n666), .C1(new_n673), .C2(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n677), .A2(new_n447), .A3(new_n476), .A4(new_n475), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT45), .Z(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n459), .B2(new_n665), .ZN(new_n681));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n664), .C1(new_n673), .C2(new_n676), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n546), .A2(new_n547), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n663), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n448), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n476), .B2(new_n475), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n679), .A2(new_n688), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n677), .A2(G36gat), .A3(new_n456), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n681), .A2(new_n669), .A3(new_n682), .A4(new_n686), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G36gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n691), .B(KEYINPUT105), .C1(new_n695), .C2(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(new_n655), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n702), .A3(new_n686), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G43gat), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n677), .A2(G43gat), .A3(new_n442), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1330gat));
  NAND3_X1  g508(.A1(new_n683), .A2(new_n446), .A3(new_n686), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n713), .A2(new_n490), .A3(new_n446), .A4(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n711), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n711), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NOR4_X1   g517(.A1(new_n684), .A2(new_n664), .A3(new_n662), .A4(new_n645), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n460), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n447), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT107), .B(G57gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n456), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  INV_X1    g527(.A(G71gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n720), .B2(new_n442), .ZN(new_n730));
  INV_X1    g529(.A(new_n720), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n655), .A2(new_n729), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n446), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n685), .A2(new_n662), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT109), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n664), .B(new_n740), .C1(new_n673), .C2(new_n676), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n645), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n745), .A2(new_n597), .A3(new_n448), .A4(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n740), .A2(new_n746), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n683), .A2(new_n448), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n597), .B2(new_n749), .ZN(G1336gat));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n456), .A2(G92gat), .A3(new_n645), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n743), .B2(new_n744), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n681), .A2(new_n669), .A3(new_n682), .A4(new_n748), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n742), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n759), .A3(KEYINPUT51), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n752), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n763), .B2(new_n755), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n751), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n741), .A2(new_n759), .A3(KEYINPUT51), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT51), .B1(new_n741), .B2(new_n759), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n768), .A2(new_n752), .B1(G92gat), .B2(new_n754), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT111), .B(new_n757), .C1(new_n769), .C2(new_n756), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n770), .ZN(G1337gat));
  NOR3_X1   g570(.A1(new_n442), .A2(G99gat), .A3(new_n645), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT113), .Z(new_n773));
  NAND2_X1  g572(.A1(new_n745), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n683), .A2(new_n702), .A3(new_n748), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G99gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n256), .A2(G106gat), .A3(new_n645), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n743), .B2(new_n744), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n681), .A2(new_n446), .A3(new_n682), .A4(new_n748), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT114), .B(G106gat), .Z(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n761), .A2(new_n762), .A3(new_n781), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n785), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n768), .A2(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n792), .B(new_n787), .C1(new_n793), .C2(new_n786), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n630), .A2(new_n632), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n624), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n607), .A2(new_n610), .A3(new_n625), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n637), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n641), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n637), .A3(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n636), .A2(new_n802), .A3(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n642), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n803), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n536), .A2(new_n537), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n525), .B1(new_n524), .B2(new_n527), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n466), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n546), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n664), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT116), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n808), .A2(new_n684), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n746), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n665), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n583), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n646), .A2(new_n685), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n675), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n447), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n684), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n549), .A2(new_n328), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n824), .B2(new_n826), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n746), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n583), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n325), .A3(new_n664), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT117), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n824), .A2(new_n835), .A3(new_n325), .A4(new_n664), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n833), .A2(KEYINPUT118), .A3(new_n834), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n325), .B1(new_n824), .B2(new_n664), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n833), .A2(new_n836), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1343gat));
  INV_X1    g644(.A(new_n205), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n446), .C1(new_n819), .C2(new_n821), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n702), .A2(new_n447), .A3(new_n669), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n813), .B(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n807), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n801), .A2(KEYINPUT119), .A3(new_n803), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n805), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n545), .B2(new_n548), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n664), .B1(new_n857), .B2(new_n816), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n662), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n820), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n847), .B1(new_n860), .B2(new_n446), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n850), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n846), .B1(new_n863), .B2(new_n549), .ZN(new_n864));
  INV_X1    g663(.A(new_n822), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n702), .A2(new_n256), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n448), .A2(new_n865), .A3(new_n456), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n218), .A3(new_n550), .ZN(new_n868));
  XOR2_X1   g667(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n846), .B1(new_n863), .B2(new_n685), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n868), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n207), .A3(new_n746), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n684), .A2(new_n461), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n546), .A2(KEYINPUT96), .A3(new_n547), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n646), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n549), .A2(KEYINPUT121), .A3(new_n646), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n636), .A2(new_n802), .A3(KEYINPUT54), .ZN(new_n884));
  INV_X1    g683(.A(new_n641), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n636), .B2(KEYINPUT54), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n853), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n806), .A3(new_n855), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n804), .A2(new_n642), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n877), .B2(new_n878), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n665), .B1(new_n891), .B2(new_n817), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n813), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(new_n662), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT122), .B(new_n847), .C1(new_n894), .C2(new_n256), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  INV_X1    g695(.A(new_n813), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n662), .B1(new_n858), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n881), .A2(new_n882), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n256), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n446), .C1(new_n819), .C2(new_n821), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n849), .A2(new_n746), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n876), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n876), .A2(G148gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n862), .B2(new_n746), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n875), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT123), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n875), .C1(new_n906), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n863), .B2(new_n662), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n867), .A2(new_n215), .A3(new_n583), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  AOI21_X1  g715(.A(G162gat), .B1(new_n867), .B2(new_n664), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n665), .A2(new_n216), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n862), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n456), .A2(new_n448), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n452), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n865), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n265), .A3(new_n549), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n822), .A2(new_n448), .A3(new_n456), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n452), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n684), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(new_n265), .ZN(G1348gat));
  OAI21_X1  g728(.A(G176gat), .B1(new_n923), .B2(new_n645), .ZN(new_n930));
  INV_X1    g729(.A(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n746), .A2(new_n266), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n923), .B2(new_n662), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n662), .A2(new_n258), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n934), .B(new_n935), .C1(new_n926), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g738(.A1(new_n665), .A2(G190gat), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n664), .A3(new_n865), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(G190gat), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n942), .A2(new_n941), .A3(G190gat), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n931), .A2(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n866), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n684), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n655), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT127), .Z(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(new_n903), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n550), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  NOR3_X1   g752(.A1(new_n946), .A2(G204gat), .A3(new_n645), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(new_n746), .A3(new_n903), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n947), .A2(new_n227), .A3(new_n583), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n949), .A2(new_n662), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n227), .B1(new_n903), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(KEYINPUT63), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  NAND2_X1  g763(.A1(new_n951), .A2(new_n664), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G218gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n228), .A3(new_n664), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


