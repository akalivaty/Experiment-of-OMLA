

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736;

  NAND2_X1 U361 ( .A1(n360), .A2(n359), .ZN(n358) );
  AND2_X1 U362 ( .A1(n649), .A2(n370), .ZN(n515) );
  XNOR2_X1 U363 ( .A(n452), .B(n714), .ZN(n442) );
  XNOR2_X1 U364 ( .A(n413), .B(G134), .ZN(n438) );
  INV_X1 U365 ( .A(KEYINPUT64), .ZN(n349) );
  INV_X1 U366 ( .A(KEYINPUT65), .ZN(n371) );
  NOR2_X1 U367 ( .A1(G953), .A2(G237), .ZN(n446) );
  NOR2_X2 U368 ( .A1(n526), .A2(KEYINPUT81), .ZN(n521) );
  NOR2_X2 U369 ( .A1(n511), .A2(n510), .ZN(n530) );
  XNOR2_X2 U370 ( .A(n398), .B(n397), .ZN(n495) );
  AND2_X2 U371 ( .A1(n574), .A2(n396), .ZN(n398) );
  NOR2_X1 U372 ( .A1(n483), .A2(n487), .ZN(n484) );
  INV_X8 U373 ( .A(G953), .ZN(n730) );
  NOR2_X1 U374 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U375 ( .A(n721), .B(n381), .ZN(n452) );
  XNOR2_X1 U376 ( .A(n348), .B(n347), .ZN(n721) );
  XNOR2_X1 U377 ( .A(n356), .B(n355), .ZN(n413) );
  XNOR2_X2 U378 ( .A(G125), .B(G140), .ZN(n418) );
  NOR2_X2 U379 ( .A1(G902), .A2(n691), .ZN(n445) );
  XNOR2_X2 U380 ( .A(n433), .B(n432), .ZN(n520) );
  NOR2_X2 U381 ( .A1(G902), .A2(n693), .ZN(n433) );
  XNOR2_X2 U382 ( .A(n454), .B(KEYINPUT85), .ZN(n722) );
  XNOR2_X2 U383 ( .A(n438), .B(n437), .ZN(n454) );
  INV_X1 U384 ( .A(n631), .ZN(n341) );
  XNOR2_X1 U385 ( .A(n387), .B(n386), .ZN(n535) );
  XNOR2_X1 U386 ( .A(n385), .B(KEYINPUT76), .ZN(n386) );
  AND2_X1 U387 ( .A1(n344), .A2(n459), .ZN(n482) );
  XNOR2_X1 U388 ( .A(n346), .B(n345), .ZN(n344) );
  INV_X1 U389 ( .A(KEYINPUT106), .ZN(n345) );
  XNOR2_X1 U390 ( .A(n560), .B(n559), .ZN(n590) );
  AND2_X1 U391 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U392 ( .A(n413), .ZN(n366) );
  INV_X1 U393 ( .A(KEYINPUT39), .ZN(n542) );
  XNOR2_X1 U394 ( .A(n518), .B(n361), .ZN(n360) );
  INV_X1 U395 ( .A(KEYINPUT34), .ZN(n361) );
  XNOR2_X1 U396 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U397 ( .A(n477), .B(n476), .ZN(n547) );
  XNOR2_X1 U398 ( .A(n475), .B(KEYINPUT25), .ZN(n476) );
  OR2_X2 U399 ( .A1(n495), .A2(n435), .ZN(n367) );
  XNOR2_X1 U400 ( .A(n547), .B(n478), .ZN(n652) );
  INV_X1 U401 ( .A(KEYINPUT104), .ZN(n478) );
  NOR2_X1 U402 ( .A1(n730), .A2(G952), .ZN(n702) );
  XNOR2_X1 U403 ( .A(n594), .B(n353), .ZN(n544) );
  INV_X1 U404 ( .A(KEYINPUT38), .ZN(n353) );
  XNOR2_X1 U405 ( .A(G146), .B(KEYINPUT67), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n349), .B(KEYINPUT4), .ZN(n348) );
  XOR2_X1 U407 ( .A(KEYINPUT7), .B(G122), .Z(n404) );
  XOR2_X1 U408 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n406) );
  XNOR2_X1 U409 ( .A(KEYINPUT10), .B(n419), .ZN(n723) );
  XNOR2_X1 U410 ( .A(KEYINPUT75), .B(G143), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n371), .B(G128), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n372), .B(KEYINPUT17), .ZN(n365) );
  NOR2_X1 U413 ( .A1(n544), .A2(n352), .ZN(n369) );
  INV_X1 U414 ( .A(n569), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n589), .B(n588), .ZN(n599) );
  XNOR2_X1 U416 ( .A(G146), .B(n723), .ZN(n466) );
  XOR2_X1 U417 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n424) );
  XNOR2_X1 U418 ( .A(n450), .B(n380), .ZN(n716) );
  XNOR2_X1 U419 ( .A(n379), .B(G122), .ZN(n380) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n736) );
  XNOR2_X1 U421 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n350) );
  NOR2_X1 U422 ( .A1(n566), .A2(n565), .ZN(n644) );
  INV_X1 U423 ( .A(KEYINPUT35), .ZN(n357) );
  INV_X1 U424 ( .A(KEYINPUT32), .ZN(n343) );
  XNOR2_X1 U425 ( .A(n480), .B(n362), .ZN(n511) );
  INV_X1 U426 ( .A(KEYINPUT105), .ZN(n362) );
  NOR2_X1 U427 ( .A1(n696), .A2(n702), .ZN(n697) );
  XNOR2_X1 U428 ( .A(n340), .B(n339), .ZN(n692) );
  XNOR2_X1 U429 ( .A(n511), .B(n381), .ZN(G3) );
  NOR2_X1 U430 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U431 ( .A1(n620), .A2(n702), .ZN(n622) );
  NOR2_X1 U432 ( .A1(n611), .A2(n702), .ZN(n613) );
  XNOR2_X1 U433 ( .A(n691), .B(n690), .ZN(n339) );
  NAND2_X1 U434 ( .A1(n698), .A2(G469), .ZN(n340) );
  NOR2_X4 U435 ( .A1(n648), .A2(n601), .ZN(n698) );
  NAND2_X1 U436 ( .A1(n342), .A2(n341), .ZN(n512) );
  XNOR2_X1 U437 ( .A(n342), .B(G119), .ZN(G21) );
  XNOR2_X1 U438 ( .A(n484), .B(n343), .ZN(n342) );
  NAND2_X1 U439 ( .A1(n649), .A2(n652), .ZN(n346) );
  XNOR2_X2 U440 ( .A(n354), .B(KEYINPUT1), .ZN(n649) );
  NOR2_X1 U441 ( .A1(n734), .A2(n736), .ZN(n554) );
  NAND2_X1 U442 ( .A1(n596), .A2(n639), .ZN(n351) );
  AND2_X1 U443 ( .A1(n354), .A2(n370), .ZN(n492) );
  XNOR2_X1 U444 ( .A(n354), .B(KEYINPUT110), .ZN(n551) );
  XNOR2_X2 U445 ( .A(n445), .B(n444), .ZN(n354) );
  INV_X1 U446 ( .A(n614), .ZN(n526) );
  XNOR2_X2 U447 ( .A(n358), .B(n357), .ZN(n614) );
  INV_X1 U448 ( .A(n573), .ZN(n359) );
  XNOR2_X1 U449 ( .A(n716), .B(n363), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n364), .B(n366), .ZN(n363) );
  XNOR2_X1 U451 ( .A(n375), .B(n365), .ZN(n364) );
  NOR2_X1 U452 ( .A1(n487), .A2(n460), .ZN(n462) );
  XNOR2_X2 U453 ( .A(n367), .B(KEYINPUT22), .ZN(n487) );
  XNOR2_X1 U454 ( .A(n603), .B(n602), .ZN(n605) );
  NAND2_X1 U455 ( .A1(n698), .A2(G478), .ZN(n603) );
  NOR2_X1 U456 ( .A1(n479), .A2(n652), .ZN(n480) );
  XOR2_X1 U457 ( .A(n469), .B(KEYINPUT89), .Z(n368) );
  AND2_X1 U458 ( .A1(n547), .A2(n490), .ZN(n370) );
  INV_X1 U459 ( .A(KEYINPUT45), .ZN(n531) );
  INV_X1 U460 ( .A(KEYINPUT107), .ZN(n559) );
  INV_X1 U461 ( .A(G469), .ZN(n444) );
  INV_X1 U462 ( .A(KEYINPUT48), .ZN(n588) );
  INV_X1 U463 ( .A(KEYINPUT16), .ZN(n379) );
  XNOR2_X1 U464 ( .A(n368), .B(n471), .ZN(n472) );
  INV_X1 U465 ( .A(n702), .ZN(n604) );
  INV_X1 U466 ( .A(KEYINPUT63), .ZN(n612) );
  INV_X1 U467 ( .A(KEYINPUT124), .ZN(n606) );
  NAND2_X1 U468 ( .A1(G224), .A2(n730), .ZN(n372) );
  XOR2_X1 U469 ( .A(KEYINPUT73), .B(KEYINPUT18), .Z(n374) );
  XNOR2_X1 U470 ( .A(G125), .B(KEYINPUT83), .ZN(n373) );
  XNOR2_X1 U471 ( .A(n374), .B(n373), .ZN(n375) );
  INV_X1 U472 ( .A(KEYINPUT3), .ZN(n376) );
  XNOR2_X1 U473 ( .A(n376), .B(G119), .ZN(n378) );
  XNOR2_X1 U474 ( .A(G116), .B(G113), .ZN(n377) );
  XNOR2_X1 U475 ( .A(n378), .B(n377), .ZN(n450) );
  INV_X1 U476 ( .A(G101), .ZN(n381) );
  XOR2_X1 U477 ( .A(G107), .B(G104), .Z(n382) );
  XNOR2_X1 U478 ( .A(G110), .B(n382), .ZN(n714) );
  XNOR2_X1 U479 ( .A(n383), .B(n442), .ZN(n615) );
  XNOR2_X1 U480 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n384) );
  XNOR2_X1 U481 ( .A(n384), .B(G902), .ZN(n601) );
  NAND2_X1 U482 ( .A1(n615), .A2(n601), .ZN(n387) );
  OR2_X1 U483 ( .A1(G902), .A2(G237), .ZN(n388) );
  NAND2_X1 U484 ( .A1(n388), .A2(G210), .ZN(n385) );
  NAND2_X1 U485 ( .A1(G214), .A2(n388), .ZN(n666) );
  INV_X1 U486 ( .A(n666), .ZN(n389) );
  NOR2_X2 U487 ( .A1(n535), .A2(n389), .ZN(n561) );
  XOR2_X1 U488 ( .A(KEYINPUT72), .B(KEYINPUT19), .Z(n390) );
  XNOR2_X1 U489 ( .A(n561), .B(n390), .ZN(n574) );
  NOR2_X1 U490 ( .A1(G898), .A2(n730), .ZN(n718) );
  NAND2_X1 U491 ( .A1(G237), .A2(G234), .ZN(n391) );
  XNOR2_X1 U492 ( .A(n391), .B(KEYINPUT14), .ZN(n393) );
  NAND2_X1 U493 ( .A1(G902), .A2(n393), .ZN(n536) );
  INV_X1 U494 ( .A(n536), .ZN(n392) );
  NAND2_X1 U495 ( .A1(n718), .A2(n392), .ZN(n395) );
  NAND2_X1 U496 ( .A1(G952), .A2(n393), .ZN(n679) );
  NOR2_X1 U497 ( .A1(G953), .A2(n679), .ZN(n394) );
  XOR2_X1 U498 ( .A(KEYINPUT84), .B(n394), .Z(n539) );
  NAND2_X1 U499 ( .A1(n395), .A2(n539), .ZN(n396) );
  INV_X1 U500 ( .A(KEYINPUT0), .ZN(n397) );
  NAND2_X1 U501 ( .A1(n601), .A2(G234), .ZN(n400) );
  XNOR2_X1 U502 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n399) );
  XNOR2_X1 U503 ( .A(n400), .B(n399), .ZN(n474) );
  NAND2_X1 U504 ( .A1(G221), .A2(n474), .ZN(n402) );
  XOR2_X1 U505 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n401) );
  XNOR2_X1 U506 ( .A(n402), .B(n401), .ZN(n653) );
  XNOR2_X1 U507 ( .A(n653), .B(KEYINPUT92), .ZN(n489) );
  XNOR2_X1 U508 ( .A(G107), .B(G116), .ZN(n403) );
  XNOR2_X1 U509 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U510 ( .A(KEYINPUT9), .B(KEYINPUT99), .ZN(n405) );
  XNOR2_X1 U511 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U512 ( .A(n408), .B(n407), .Z(n412) );
  XOR2_X1 U513 ( .A(KEYINPUT78), .B(KEYINPUT8), .Z(n410) );
  NAND2_X1 U514 ( .A1(G234), .A2(n730), .ZN(n409) );
  XNOR2_X1 U515 ( .A(n410), .B(n409), .ZN(n470) );
  NAND2_X1 U516 ( .A1(G217), .A2(n470), .ZN(n411) );
  XNOR2_X1 U517 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U518 ( .A(n414), .B(n438), .ZN(n602) );
  INV_X1 U519 ( .A(G902), .ZN(n415) );
  NAND2_X1 U520 ( .A1(n602), .A2(n415), .ZN(n417) );
  XOR2_X1 U521 ( .A(G478), .B(KEYINPUT101), .Z(n416) );
  XNOR2_X1 U522 ( .A(n417), .B(n416), .ZN(n519) );
  INV_X1 U523 ( .A(n519), .ZN(n498) );
  INV_X1 U524 ( .A(n418), .ZN(n419) );
  XOR2_X1 U525 ( .A(KEYINPUT11), .B(G113), .Z(n421) );
  XNOR2_X1 U526 ( .A(G143), .B(G122), .ZN(n420) );
  XNOR2_X1 U527 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U528 ( .A(n466), .B(n422), .ZN(n429) );
  NAND2_X1 U529 ( .A1(n446), .A2(G214), .ZN(n423) );
  XNOR2_X1 U530 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U531 ( .A(n425), .B(KEYINPUT12), .Z(n427) );
  XNOR2_X1 U532 ( .A(G104), .B(G131), .ZN(n426) );
  XNOR2_X1 U533 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U534 ( .A(n429), .B(n428), .ZN(n693) );
  XNOR2_X1 U535 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n431) );
  INV_X1 U536 ( .A(G475), .ZN(n430) );
  INV_X1 U537 ( .A(n520), .ZN(n499) );
  NAND2_X1 U538 ( .A1(n498), .A2(n499), .ZN(n668) );
  NOR2_X1 U539 ( .A1(n489), .A2(n668), .ZN(n434) );
  XNOR2_X1 U540 ( .A(n434), .B(KEYINPUT103), .ZN(n435) );
  XNOR2_X1 U541 ( .A(G137), .B(G131), .ZN(n436) );
  XNOR2_X1 U542 ( .A(n436), .B(KEYINPUT68), .ZN(n437) );
  XOR2_X1 U543 ( .A(KEYINPUT86), .B(G140), .Z(n440) );
  NAND2_X1 U544 ( .A1(G227), .A2(n730), .ZN(n439) );
  XNOR2_X1 U545 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U547 ( .A(n722), .B(n443), .ZN(n691) );
  INV_X1 U548 ( .A(n649), .ZN(n566) );
  NAND2_X1 U549 ( .A1(n446), .A2(G210), .ZN(n447) );
  XNOR2_X1 U550 ( .A(n447), .B(KEYINPUT71), .ZN(n449) );
  XNOR2_X1 U551 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n448) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U555 ( .A(n454), .B(n455), .ZN(n608) );
  OR2_X1 U556 ( .A1(n608), .A2(G902), .ZN(n458) );
  INV_X1 U557 ( .A(KEYINPUT70), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n456), .B(G472), .ZN(n457) );
  XNOR2_X2 U559 ( .A(n458), .B(n457), .ZN(n549) );
  XNOR2_X1 U560 ( .A(n549), .B(KEYINPUT6), .ZN(n557) );
  INV_X1 U561 ( .A(n557), .ZN(n459) );
  NAND2_X1 U562 ( .A1(n566), .A2(n459), .ZN(n460) );
  INV_X1 U563 ( .A(KEYINPUT80), .ZN(n461) );
  XNOR2_X1 U564 ( .A(n462), .B(n461), .ZN(n479) );
  XOR2_X1 U565 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n464) );
  XNOR2_X1 U566 ( .A(G128), .B(G137), .ZN(n463) );
  XNOR2_X1 U567 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n466), .B(n465), .ZN(n473) );
  XOR2_X1 U569 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n468) );
  XNOR2_X1 U570 ( .A(G110), .B(G119), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U572 ( .A1(G221), .A2(n470), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n473), .B(n472), .ZN(n699) );
  NOR2_X1 U574 ( .A1(G902), .A2(n699), .ZN(n477) );
  NAND2_X1 U575 ( .A1(G217), .A2(n474), .ZN(n475) );
  INV_X1 U576 ( .A(KEYINPUT74), .ZN(n481) );
  XNOR2_X1 U577 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U578 ( .A(n549), .ZN(n658) );
  NOR2_X1 U579 ( .A1(n547), .A2(n658), .ZN(n485) );
  NAND2_X1 U580 ( .A1(n566), .A2(n485), .ZN(n486) );
  NOR2_X1 U581 ( .A1(n487), .A2(n486), .ZN(n631) );
  NOR2_X1 U582 ( .A1(KEYINPUT44), .A2(KEYINPUT69), .ZN(n513) );
  INV_X1 U583 ( .A(n513), .ZN(n488) );
  NAND2_X1 U584 ( .A1(n512), .A2(n488), .ZN(n509) );
  INV_X1 U585 ( .A(n495), .ZN(n517) );
  INV_X1 U586 ( .A(n489), .ZN(n490) );
  AND2_X1 U587 ( .A1(n515), .A2(n658), .ZN(n661) );
  NAND2_X1 U588 ( .A1(n517), .A2(n661), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n491), .B(KEYINPUT31), .ZN(n642) );
  INV_X1 U590 ( .A(n642), .ZN(n497) );
  XNOR2_X1 U591 ( .A(n492), .B(KEYINPUT93), .ZN(n567) );
  INV_X1 U592 ( .A(n567), .ZN(n493) );
  NAND2_X1 U593 ( .A1(n493), .A2(n549), .ZN(n494) );
  NOR2_X1 U594 ( .A1(n495), .A2(n494), .ZN(n626) );
  INV_X1 U595 ( .A(n626), .ZN(n496) );
  NAND2_X1 U596 ( .A1(n497), .A2(n496), .ZN(n501) );
  NOR2_X1 U597 ( .A1(n498), .A2(n520), .ZN(n641) );
  NOR2_X4 U598 ( .A1(n499), .A2(n519), .ZN(n639) );
  OR2_X1 U599 ( .A1(n641), .A2(n639), .ZN(n500) );
  XNOR2_X1 U600 ( .A(KEYINPUT102), .B(n500), .ZN(n669) );
  XOR2_X1 U601 ( .A(KEYINPUT77), .B(n669), .Z(n577) );
  NAND2_X1 U602 ( .A1(n501), .A2(n577), .ZN(n507) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n523) );
  INV_X1 U604 ( .A(KEYINPUT81), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n523), .A2(n502), .ZN(n505) );
  INV_X1 U606 ( .A(KEYINPUT69), .ZN(n503) );
  NAND2_X1 U607 ( .A1(n503), .A2(KEYINPUT44), .ZN(n504) );
  NAND2_X1 U608 ( .A1(n505), .A2(n504), .ZN(n506) );
  AND2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U610 ( .A1(n509), .A2(n508), .ZN(n510) );
  INV_X1 U611 ( .A(n512), .ZN(n514) );
  NAND2_X1 U612 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U613 ( .A1(n515), .A2(n557), .ZN(n516) );
  XNOR2_X2 U614 ( .A(n516), .B(KEYINPUT33), .ZN(n683) );
  NAND2_X1 U615 ( .A1(n683), .A2(n517), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n520), .A2(n519), .ZN(n573) );
  NAND2_X1 U617 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U618 ( .A1(n523), .A2(KEYINPUT81), .ZN(n524) );
  NOR2_X1 U619 ( .A1(n524), .A2(KEYINPUT69), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U622 ( .A1(n529), .A2(n530), .ZN(n532) );
  XNOR2_X2 U623 ( .A(n532), .B(n531), .ZN(n709) );
  NAND2_X1 U624 ( .A1(n658), .A2(n666), .ZN(n534) );
  XOR2_X1 U625 ( .A(KEYINPUT30), .B(KEYINPUT109), .Z(n533) );
  XNOR2_X1 U626 ( .A(n534), .B(n533), .ZN(n568) );
  INV_X1 U627 ( .A(n568), .ZN(n540) );
  BUF_X1 U628 ( .A(n535), .Z(n594) );
  NOR2_X1 U629 ( .A1(G900), .A2(n536), .ZN(n537) );
  NAND2_X1 U630 ( .A1(G953), .A2(n537), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n540), .A2(n369), .ZN(n541) );
  NOR2_X1 U633 ( .A1(n567), .A2(n541), .ZN(n543) );
  XNOR2_X1 U634 ( .A(n543), .B(n542), .ZN(n596) );
  INV_X1 U635 ( .A(n544), .ZN(n665) );
  NAND2_X1 U636 ( .A1(n666), .A2(n665), .ZN(n671) );
  NOR2_X1 U637 ( .A1(n671), .A2(n668), .ZN(n546) );
  XNOR2_X1 U638 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n681) );
  NOR2_X1 U640 ( .A1(n653), .A2(n547), .ZN(n548) );
  NAND2_X1 U641 ( .A1(n548), .A2(n569), .ZN(n555) );
  NOR2_X1 U642 ( .A1(n555), .A2(n549), .ZN(n550) );
  XNOR2_X1 U643 ( .A(n550), .B(KEYINPUT28), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n575) );
  NOR2_X1 U645 ( .A1(n681), .A2(n575), .ZN(n553) );
  XNOR2_X1 U646 ( .A(KEYINPUT42), .B(n553), .ZN(n734) );
  XNOR2_X1 U647 ( .A(n554), .B(KEYINPUT46), .ZN(n587) );
  INV_X1 U648 ( .A(n639), .ZN(n556) );
  NOR2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U650 ( .A(n590), .ZN(n563) );
  INV_X1 U651 ( .A(n561), .ZN(n562) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(n564), .Z(n565) );
  XNOR2_X1 U653 ( .A(KEYINPUT79), .B(n644), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U655 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U656 ( .A1(n571), .A2(n594), .ZN(n572) );
  NOR2_X1 U657 ( .A1(n573), .A2(n572), .ZN(n634) );
  XNOR2_X1 U658 ( .A(KEYINPUT47), .B(KEYINPUT66), .ZN(n579) );
  INV_X1 U659 ( .A(n574), .ZN(n576) );
  NOR2_X1 U660 ( .A1(n576), .A2(n575), .ZN(n636) );
  NAND2_X1 U661 ( .A1(n636), .A2(n577), .ZN(n578) );
  NOR2_X1 U662 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U663 ( .A1(n634), .A2(n580), .ZN(n581) );
  NAND2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n636), .A2(n669), .ZN(n583) );
  AND2_X1 U666 ( .A1(n583), .A2(KEYINPUT47), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n666), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n649), .A2(n591), .ZN(n593) );
  XOR2_X1 U670 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n592) );
  XNOR2_X1 U671 ( .A(n593), .B(n592), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n647) );
  AND2_X1 U673 ( .A1(n596), .A2(n641), .ZN(n646) );
  INV_X1 U674 ( .A(n646), .ZN(n597) );
  AND2_X1 U675 ( .A1(n647), .A2(n597), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n728) );
  NOR2_X2 U677 ( .A1(n709), .A2(n728), .ZN(n600) );
  XNOR2_X2 U678 ( .A(n600), .B(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(n606), .ZN(G63) );
  NAND2_X1 U681 ( .A1(n698), .A2(G472), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT62), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n613), .B(n612), .ZN(G57) );
  XNOR2_X1 U685 ( .A(n614), .B(G122), .ZN(G24) );
  NAND2_X1 U686 ( .A1(n698), .A2(G210), .ZN(n619) );
  XNOR2_X1 U687 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n616), .B(KEYINPUT55), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n615), .B(n617), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  XOR2_X1 U691 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G51) );
  NAND2_X1 U693 ( .A1(n626), .A2(n639), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(G104), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n625) );
  XNOR2_X1 U696 ( .A(KEYINPUT26), .B(KEYINPUT27), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n630) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT113), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n641), .A2(n626), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(G9) );
  XOR2_X1 U702 ( .A(G110), .B(n631), .Z(G12) );
  XOR2_X1 U703 ( .A(G128), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U704 ( .A1(n636), .A2(n641), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(G30) );
  XOR2_X1 U706 ( .A(G143), .B(n634), .Z(n635) );
  XNOR2_X1 U707 ( .A(KEYINPUT116), .B(n635), .ZN(G45) );
  XOR2_X1 U708 ( .A(G146), .B(KEYINPUT117), .Z(n638) );
  NAND2_X1 U709 ( .A1(n636), .A2(n639), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n642), .A2(n639), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(G113), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(G116), .ZN(G18) );
  XNOR2_X1 U715 ( .A(G125), .B(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U717 ( .A(G134), .B(n646), .Z(G36) );
  XNOR2_X1 U718 ( .A(G140), .B(n647), .ZN(G42) );
  INV_X1 U719 ( .A(n648), .ZN(n687) );
  NOR2_X1 U720 ( .A1(n370), .A2(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n657) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n655) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT120), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT51), .B(n663), .Z(n664) );
  NOR2_X1 U731 ( .A1(n681), .A2(n664), .ZN(n676) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n673) );
  INV_X1 U734 ( .A(n669), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  AND2_X1 U737 ( .A1(n683), .A2(n674), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT121), .ZN(n685) );
  INV_X1 U742 ( .A(n681), .ZN(n682) );
  NAND2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U746 ( .A1(n730), .A2(n688), .ZN(n689) );
  XOR2_X1 U747 ( .A(KEYINPUT53), .B(n689), .Z(G75) );
  XOR2_X1 U748 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n690) );
  NOR2_X1 U749 ( .A1(n702), .A2(n692), .ZN(G54) );
  NAND2_X1 U750 ( .A1(n698), .A2(G475), .ZN(n695) );
  XOR2_X1 U751 ( .A(n693), .B(KEYINPUT59), .Z(n694) );
  XNOR2_X1 U752 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n697), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n698), .A2(G217), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U756 ( .A1(n702), .A2(n701), .ZN(G66) );
  NAND2_X1 U757 ( .A1(G224), .A2(KEYINPUT61), .ZN(n707) );
  INV_X1 U758 ( .A(G898), .ZN(n705) );
  AND2_X1 U759 ( .A1(G953), .A2(G224), .ZN(n703) );
  NOR2_X1 U760 ( .A1(KEYINPUT61), .A2(n703), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U763 ( .A1(G898), .A2(KEYINPUT61), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U765 ( .A1(n710), .A2(n730), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n713), .B(KEYINPUT125), .ZN(n720) );
  XOR2_X1 U768 ( .A(G101), .B(n714), .Z(n715) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U771 ( .A(n720), .B(n719), .Z(G69) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n729) );
  XNOR2_X1 U774 ( .A(n729), .B(KEYINPUT126), .ZN(n725) );
  XNOR2_X1 U775 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U776 ( .A1(G900), .A2(n726), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G953), .ZN(n733) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U781 ( .A(G137), .B(KEYINPUT127), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(G39) );
  XOR2_X1 U783 ( .A(G131), .B(n736), .Z(G33) );
endmodule

