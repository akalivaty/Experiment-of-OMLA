

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776;

  XOR2_X1 U370 ( .A(n691), .B(n690), .Z(n357) );
  XOR2_X1 U371 ( .A(n680), .B(KEYINPUT121), .Z(n361) );
  XOR2_X1 U372 ( .A(n683), .B(n682), .Z(n360) );
  AND2_X1 U373 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X1 U374 ( .A1(n446), .A2(n444), .ZN(n454) );
  NOR2_X1 U375 ( .A1(n400), .A2(n352), .ZN(n670) );
  BUF_X1 U376 ( .A(n599), .Z(n347) );
  OR2_X1 U377 ( .A1(n408), .A2(n627), .ZN(n401) );
  NOR2_X1 U378 ( .A1(n625), .A2(n666), .ZN(n644) );
  AND2_X1 U379 ( .A1(n586), .A2(n423), .ZN(n624) );
  XNOR2_X1 U380 ( .A(n754), .B(n522), .ZN(n691) );
  XNOR2_X1 U381 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n496) );
  XNOR2_X1 U382 ( .A(G113), .B(G101), .ZN(n498) );
  NAND2_X1 U383 ( .A1(n375), .A2(n376), .ZN(n594) );
  XNOR2_X2 U384 ( .A(n626), .B(KEYINPUT19), .ZN(n532) );
  XNOR2_X1 U385 ( .A(n598), .B(KEYINPUT106), .ZN(n634) );
  AND2_X4 U386 ( .A1(n368), .A2(n367), .ZN(n689) );
  XNOR2_X2 U387 ( .A(n505), .B(KEYINPUT95), .ZN(n765) );
  AND2_X2 U388 ( .A1(n378), .A2(n377), .ZN(n376) );
  XOR2_X1 U389 ( .A(KEYINPUT4), .B(G146), .Z(n515) );
  XNOR2_X1 U390 ( .A(G110), .B(G128), .ZN(n473) );
  INV_X2 U391 ( .A(G953), .ZN(n767) );
  AND2_X2 U392 ( .A1(n433), .A2(n432), .ZN(n431) );
  AND2_X2 U393 ( .A1(n365), .A2(n380), .ZN(n355) );
  AND2_X1 U394 ( .A1(n452), .A2(n451), .ZN(n378) );
  INV_X1 U395 ( .A(n724), .ZN(n453) );
  NOR2_X1 U396 ( .A1(n713), .A2(n616), .ZN(n369) );
  OR2_X1 U397 ( .A1(n706), .A2(n374), .ZN(n371) );
  XNOR2_X1 U398 ( .A(n629), .B(KEYINPUT82), .ZN(n706) );
  AND2_X1 U399 ( .A1(n373), .A2(n661), .ZN(n372) );
  OR2_X1 U400 ( .A1(n630), .A2(n374), .ZN(n373) );
  OR2_X1 U401 ( .A1(n580), .A2(n581), .ZN(n696) );
  NAND2_X1 U402 ( .A1(n618), .A2(n495), .ZN(n710) );
  XNOR2_X2 U403 ( .A(n348), .B(n349), .ZN(n615) );
  NOR2_X1 U404 ( .A1(n685), .A2(G902), .ZN(n348) );
  XOR2_X1 U405 ( .A(n470), .B(G469), .Z(n349) );
  XNOR2_X2 U406 ( .A(n350), .B(G472), .ZN(n599) );
  NOR2_X1 U407 ( .A1(n657), .A2(G902), .ZN(n350) );
  AND2_X1 U408 ( .A1(n438), .A2(n351), .ZN(n436) );
  XNOR2_X2 U409 ( .A(n611), .B(KEYINPUT39), .ZN(n649) );
  XNOR2_X2 U410 ( .A(n579), .B(n578), .ZN(n598) );
  OR2_X1 U411 ( .A1(n618), .A2(n617), .ZN(n623) );
  XNOR2_X1 U412 ( .A(n369), .B(KEYINPUT69), .ZN(n617) );
  XNOR2_X1 U413 ( .A(n640), .B(n426), .ZN(n425) );
  INV_X1 U414 ( .A(KEYINPUT84), .ZN(n426) );
  INV_X1 U415 ( .A(n623), .ZN(n423) );
  NAND2_X1 U416 ( .A1(n706), .A2(n630), .ZN(n632) );
  NOR2_X1 U417 ( .A1(n668), .A2(KEYINPUT100), .ZN(n416) );
  NOR2_X1 U418 ( .A1(n662), .A2(n460), .ZN(n442) );
  NAND2_X1 U419 ( .A1(n457), .A2(n643), .ZN(n438) );
  AND2_X1 U420 ( .A1(n665), .A2(n775), .ZN(n375) );
  NAND2_X1 U421 ( .A1(n635), .A2(n725), .ZN(n626) );
  INV_X1 U422 ( .A(KEYINPUT99), .ZN(n578) );
  XNOR2_X1 U423 ( .A(n615), .B(KEYINPUT1), .ZN(n565) );
  XNOR2_X1 U424 ( .A(G101), .B(G140), .ZN(n465) );
  INV_X1 U425 ( .A(n626), .ZN(n407) );
  NOR2_X1 U426 ( .A1(n711), .A2(n405), .ZN(n404) );
  NOR2_X1 U427 ( .A1(n407), .A2(n627), .ZN(n405) );
  NOR2_X1 U428 ( .A1(n599), .A2(n623), .ZN(n619) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n374) );
  NOR2_X1 U430 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U431 ( .A1(n663), .A2(n440), .ZN(n439) );
  NOR2_X1 U432 ( .A1(n461), .A2(KEYINPUT87), .ZN(n440) );
  NOR2_X1 U433 ( .A1(n436), .A2(n434), .ZN(n430) );
  XNOR2_X1 U434 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n549) );
  XNOR2_X1 U436 ( .A(n597), .B(KEYINPUT45), .ZN(n743) );
  XOR2_X1 U437 ( .A(G107), .B(KEYINPUT9), .Z(n539) );
  XOR2_X1 U438 ( .A(G104), .B(G122), .Z(n548) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n527) );
  INV_X1 U440 ( .A(G237), .ZN(n523) );
  INV_X1 U441 ( .A(n485), .ZN(n654) );
  INV_X1 U442 ( .A(G902), .ZN(n557) );
  XNOR2_X1 U443 ( .A(n370), .B(KEYINPUT21), .ZN(n713) );
  XNOR2_X1 U444 ( .A(n554), .B(n463), .ZN(n455) );
  XNOR2_X1 U445 ( .A(G137), .B(KEYINPUT4), .ZN(n463) );
  XNOR2_X1 U446 ( .A(G110), .B(G107), .ZN(n467) );
  BUF_X1 U447 ( .A(n743), .Z(n757) );
  NAND2_X1 U448 ( .A1(n383), .A2(n381), .ZN(n380) );
  NAND2_X1 U449 ( .A1(n654), .A2(n382), .ZN(n381) );
  OR2_X1 U450 ( .A1(n654), .A2(n655), .ZN(n383) );
  NAND2_X1 U451 ( .A1(KEYINPUT64), .A2(KEYINPUT2), .ZN(n382) );
  AND2_X1 U452 ( .A1(n654), .A2(KEYINPUT64), .ZN(n379) );
  NAND2_X1 U453 ( .A1(n366), .A2(n757), .ZN(n367) );
  AND2_X1 U454 ( .A1(n656), .A2(KEYINPUT2), .ZN(n366) );
  XNOR2_X1 U455 ( .A(G137), .B(KEYINPUT96), .ZN(n480) );
  XNOR2_X1 U456 ( .A(G119), .B(KEYINPUT23), .ZN(n481) );
  XNOR2_X1 U457 ( .A(KEYINPUT79), .B(KEYINPUT24), .ZN(n474) );
  INV_X1 U458 ( .A(G125), .ZN(n478) );
  XNOR2_X1 U459 ( .A(KEYINPUT10), .B(G140), .ZN(n479) );
  INV_X1 U460 ( .A(n367), .ZN(n745) );
  NOR2_X1 U461 ( .A1(n445), .A2(n637), .ZN(n444) );
  NOR2_X1 U462 ( .A1(n535), .A2(n536), .ZN(n445) );
  NAND2_X1 U463 ( .A1(n401), .A2(n404), .ZN(n400) );
  NOR2_X1 U464 ( .A1(n628), .A2(n421), .ZN(n629) );
  NAND2_X1 U465 ( .A1(n573), .A2(n714), .ZN(n665) );
  INV_X1 U466 ( .A(KEYINPUT122), .ZN(n386) );
  INV_X1 U467 ( .A(KEYINPUT60), .ZN(n388) );
  INV_X1 U468 ( .A(KEYINPUT120), .ZN(n390) );
  INV_X1 U469 ( .A(KEYINPUT56), .ZN(n396) );
  AND2_X1 U470 ( .A1(n441), .A2(n460), .ZN(n351) );
  INV_X1 U471 ( .A(n662), .ZN(n461) );
  AND2_X1 U472 ( .A1(n408), .A2(n406), .ZN(n352) );
  NAND2_X1 U473 ( .A1(n606), .A2(n531), .ZN(n353) );
  AND2_X1 U474 ( .A1(n535), .A2(n536), .ZN(n354) );
  XNOR2_X1 U475 ( .A(n599), .B(n506), .ZN(n586) );
  AND2_X1 U476 ( .A1(KEYINPUT34), .A2(KEYINPUT35), .ZN(n356) );
  INV_X1 U477 ( .A(KEYINPUT100), .ZN(n419) );
  XNOR2_X1 U478 ( .A(KEYINPUT88), .B(KEYINPUT46), .ZN(n358) );
  XOR2_X1 U479 ( .A(n657), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U480 ( .A(n685), .B(n687), .Z(n362) );
  INV_X1 U481 ( .A(KEYINPUT87), .ZN(n460) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(n659), .Z(n693) );
  INV_X1 U483 ( .A(n693), .ZN(n398) );
  NAND2_X1 U484 ( .A1(n355), .A2(n363), .ZN(n368) );
  NAND2_X1 U485 ( .A1(n364), .A2(n379), .ZN(n363) );
  INV_X1 U486 ( .A(n410), .ZN(n364) );
  NAND2_X1 U487 ( .A1(n410), .A2(n384), .ZN(n365) );
  NAND2_X1 U488 ( .A1(n494), .A2(G221), .ZN(n370) );
  NAND2_X1 U489 ( .A1(n372), .A2(n371), .ZN(n640) );
  NAND2_X1 U490 ( .A1(n447), .A2(n450), .ZN(n377) );
  NAND2_X1 U491 ( .A1(n377), .A2(n378), .ZN(n675) );
  AND2_X1 U492 ( .A1(n653), .A2(n655), .ZN(n384) );
  XNOR2_X1 U493 ( .A(n385), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U494 ( .A1(n392), .A2(n398), .ZN(n385) );
  XNOR2_X1 U495 ( .A(n387), .B(n386), .ZN(G63) );
  NAND2_X1 U496 ( .A1(n393), .A2(n398), .ZN(n387) );
  XNOR2_X1 U497 ( .A(n389), .B(n388), .ZN(G60) );
  NAND2_X1 U498 ( .A1(n394), .A2(n398), .ZN(n389) );
  XNOR2_X1 U499 ( .A(n391), .B(n390), .ZN(G54) );
  NAND2_X1 U500 ( .A1(n395), .A2(n398), .ZN(n391) );
  XNOR2_X1 U501 ( .A(n658), .B(n359), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n681), .B(n361), .ZN(n393) );
  XNOR2_X1 U503 ( .A(n684), .B(n360), .ZN(n394) );
  XNOR2_X1 U504 ( .A(n688), .B(n362), .ZN(n395) );
  XNOR2_X1 U505 ( .A(n397), .B(n396), .ZN(G51) );
  NAND2_X1 U506 ( .A1(n399), .A2(n398), .ZN(n397) );
  XNOR2_X1 U507 ( .A(n692), .B(n357), .ZN(n399) );
  AND2_X1 U508 ( .A1(n407), .A2(n627), .ZN(n406) );
  XNOR2_X1 U509 ( .A(n644), .B(n409), .ZN(n408) );
  INV_X1 U510 ( .A(KEYINPUT111), .ZN(n409) );
  NAND2_X1 U511 ( .A1(n652), .A2(n743), .ZN(n410) );
  NAND2_X1 U512 ( .A1(n411), .A2(n434), .ZN(n433) );
  NAND2_X1 U513 ( .A1(n437), .A2(n439), .ZN(n411) );
  INV_X1 U514 ( .A(n411), .ZN(n429) );
  AND2_X1 U515 ( .A1(n429), .A2(n412), .ZN(n656) );
  INV_X1 U516 ( .A(n436), .ZN(n412) );
  NAND2_X1 U517 ( .A1(n414), .A2(n413), .ZN(n585) );
  NAND2_X1 U518 ( .A1(n417), .A2(n668), .ZN(n413) );
  NAND2_X1 U519 ( .A1(n418), .A2(n630), .ZN(n415) );
  AND2_X1 U520 ( .A1(n696), .A2(KEYINPUT100), .ZN(n417) );
  NAND2_X1 U521 ( .A1(n420), .A2(n419), .ZN(n418) );
  INV_X1 U522 ( .A(n696), .ZN(n420) );
  XNOR2_X2 U523 ( .A(n577), .B(n576), .ZN(n668) );
  INV_X1 U524 ( .A(n532), .ZN(n421) );
  XNOR2_X2 U525 ( .A(n422), .B(KEYINPUT74), .ZN(n575) );
  NOR2_X2 U526 ( .A1(n565), .A2(n710), .ZN(n422) );
  NAND2_X1 U527 ( .A1(n427), .A2(n458), .ZN(n457) );
  XNOR2_X1 U528 ( .A(n622), .B(n358), .ZN(n427) );
  NAND2_X1 U529 ( .A1(n424), .A2(n620), .ZN(n628) );
  XNOR2_X1 U530 ( .A(n619), .B(KEYINPUT28), .ZN(n424) );
  NAND2_X1 U531 ( .A1(n641), .A2(n425), .ZN(n642) );
  NAND2_X1 U532 ( .A1(n575), .A2(n462), .ZN(n577) );
  XNOR2_X2 U533 ( .A(n443), .B(G143), .ZN(n517) );
  OR2_X2 U534 ( .A1(n574), .A2(n562), .ZN(n564) );
  NAND2_X1 U535 ( .A1(n459), .A2(n427), .ZN(n441) );
  NAND2_X1 U536 ( .A1(n431), .A2(n428), .ZN(n652) );
  NAND2_X1 U537 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U538 ( .A1(n436), .A2(n434), .ZN(n432) );
  INV_X1 U539 ( .A(KEYINPUT76), .ZN(n434) );
  NAND2_X1 U540 ( .A1(n435), .A2(n442), .ZN(n437) );
  NAND2_X1 U541 ( .A1(n438), .A2(n441), .ZN(n435) );
  XNOR2_X2 U542 ( .A(n564), .B(n563), .ZN(n589) );
  XNOR2_X2 U543 ( .A(G128), .B(KEYINPUT83), .ZN(n443) );
  NAND2_X1 U544 ( .A1(n575), .A2(n586), .ZN(n509) );
  XNOR2_X1 U545 ( .A(n575), .B(KEYINPUT51), .ZN(n709) );
  NAND2_X1 U546 ( .A1(n354), .A2(n724), .ZN(n446) );
  INV_X1 U547 ( .A(KEYINPUT35), .ZN(n448) );
  NAND2_X1 U548 ( .A1(n453), .A2(KEYINPUT34), .ZN(n449) );
  INV_X1 U549 ( .A(n454), .ZN(n450) );
  NAND2_X1 U550 ( .A1(n453), .A2(n356), .ZN(n451) );
  NAND2_X1 U551 ( .A1(n454), .A2(KEYINPUT35), .ZN(n452) );
  XNOR2_X2 U552 ( .A(n541), .B(n455), .ZN(n505) );
  XNOR2_X2 U553 ( .A(n456), .B(G131), .ZN(n554) );
  XNOR2_X2 U554 ( .A(G146), .B(KEYINPUT67), .ZN(n456) );
  XNOR2_X2 U555 ( .A(n517), .B(G134), .ZN(n541) );
  INV_X1 U556 ( .A(n642), .ZN(n458) );
  NOR2_X1 U557 ( .A1(n642), .A2(n643), .ZN(n459) );
  NOR2_X1 U558 ( .A1(n574), .A2(n347), .ZN(n462) );
  XNOR2_X1 U559 ( .A(n613), .B(n612), .ZN(n673) );
  NAND2_X1 U560 ( .A1(n767), .A2(G227), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n464), .B(KEYINPUT80), .ZN(n466) );
  XNOR2_X1 U562 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n467), .B(G104), .ZN(n511) );
  XNOR2_X1 U564 ( .A(n468), .B(n511), .ZN(n469) );
  XNOR2_X1 U565 ( .A(n765), .B(n469), .ZN(n685) );
  INV_X1 U566 ( .A(KEYINPUT70), .ZN(n470) );
  NAND2_X1 U567 ( .A1(n767), .A2(G234), .ZN(n472) );
  XNOR2_X1 U568 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n472), .B(n471), .ZN(n537) );
  NAND2_X1 U570 ( .A1(n537), .A2(G221), .ZN(n477) );
  XNOR2_X1 U571 ( .A(n473), .B(G146), .ZN(n475) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n477), .B(n476), .ZN(n484) );
  XNOR2_X1 U574 ( .A(n479), .B(n478), .ZN(n766) );
  XNOR2_X1 U575 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n766), .B(n482), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n484), .B(n483), .ZN(n676) );
  OR2_X1 U578 ( .A1(n676), .A2(G902), .ZN(n493) );
  NAND2_X1 U579 ( .A1(n485), .A2(G234), .ZN(n487) );
  XNOR2_X1 U580 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n486) );
  XNOR2_X1 U581 ( .A(n487), .B(n486), .ZN(n494) );
  AND2_X1 U582 ( .A1(n494), .A2(G217), .ZN(n491) );
  XNOR2_X1 U583 ( .A(KEYINPUT78), .B(KEYINPUT97), .ZN(n489) );
  XNOR2_X1 U584 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n488) );
  XNOR2_X1 U585 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U586 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X2 U587 ( .A(n493), .B(n492), .ZN(n618) );
  INV_X1 U588 ( .A(n713), .ZN(n495) );
  XNOR2_X1 U589 ( .A(G119), .B(G116), .ZN(n497) );
  XNOR2_X1 U590 ( .A(n497), .B(n496), .ZN(n500) );
  XNOR2_X1 U591 ( .A(n498), .B(KEYINPUT3), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n500), .B(n499), .ZN(n513) );
  XNOR2_X1 U593 ( .A(KEYINPUT75), .B(KEYINPUT5), .ZN(n502) );
  NAND2_X1 U594 ( .A1(G210), .A2(n549), .ZN(n501) );
  XNOR2_X1 U595 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n513), .B(n503), .ZN(n504) );
  XNOR2_X1 U597 ( .A(n505), .B(n504), .ZN(n657) );
  XNOR2_X1 U598 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n506) );
  XNOR2_X1 U599 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n507), .B(KEYINPUT91), .ZN(n508) );
  XNOR2_X2 U601 ( .A(n509), .B(n508), .ZN(n724) );
  XNOR2_X1 U602 ( .A(KEYINPUT16), .B(G122), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n513), .B(n512), .ZN(n754) );
  NAND2_X1 U605 ( .A1(G224), .A2(n767), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U607 ( .A(n517), .B(n516), .ZN(n521) );
  XOR2_X1 U608 ( .A(KEYINPUT18), .B(KEYINPUT92), .Z(n519) );
  XNOR2_X1 U609 ( .A(G125), .B(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U611 ( .A(n521), .B(n520), .ZN(n522) );
  OR2_X2 U612 ( .A1(n691), .A2(n654), .ZN(n525) );
  NAND2_X1 U613 ( .A1(n557), .A2(n523), .ZN(n526) );
  AND2_X1 U614 ( .A1(n526), .A2(G210), .ZN(n524) );
  XNOR2_X2 U615 ( .A(n525), .B(n524), .ZN(n635) );
  NAND2_X1 U616 ( .A1(n526), .A2(G214), .ZN(n725) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT14), .ZN(n528) );
  NAND2_X1 U618 ( .A1(G952), .A2(n528), .ZN(n738) );
  OR2_X1 U619 ( .A1(n738), .A2(G953), .ZN(n606) );
  NAND2_X1 U620 ( .A1(G902), .A2(n528), .ZN(n603) );
  INV_X1 U621 ( .A(n603), .ZN(n529) );
  NOR2_X1 U622 ( .A1(G898), .A2(n767), .ZN(n755) );
  NAND2_X1 U623 ( .A1(n529), .A2(n755), .ZN(n530) );
  XNOR2_X1 U624 ( .A(n530), .B(KEYINPUT94), .ZN(n531) );
  NAND2_X1 U625 ( .A1(n532), .A2(n353), .ZN(n534) );
  XNOR2_X1 U626 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n534), .B(n533), .ZN(n574) );
  BUF_X1 U628 ( .A(n574), .Z(n580) );
  INV_X1 U629 ( .A(n580), .ZN(n535) );
  INV_X1 U630 ( .A(KEYINPUT34), .ZN(n536) );
  NAND2_X1 U631 ( .A1(G217), .A2(n537), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U633 ( .A(n540), .B(KEYINPUT7), .Z(n544) );
  XNOR2_X1 U634 ( .A(G116), .B(G122), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n541), .B(n542), .ZN(n543) );
  XNOR2_X1 U636 ( .A(n544), .B(n543), .ZN(n680) );
  NAND2_X1 U637 ( .A1(n680), .A2(n557), .ZN(n546) );
  INV_X1 U638 ( .A(G478), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n583) );
  INV_X1 U640 ( .A(n583), .ZN(n560) );
  XNOR2_X1 U641 ( .A(G113), .B(G143), .ZN(n547) );
  XNOR2_X1 U642 ( .A(n548), .B(n547), .ZN(n553) );
  XOR2_X1 U643 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n551) );
  NAND2_X1 U644 ( .A1(G214), .A2(n549), .ZN(n550) );
  XNOR2_X1 U645 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n553), .B(n552), .ZN(n556) );
  XNOR2_X1 U647 ( .A(n554), .B(n766), .ZN(n555) );
  XNOR2_X1 U648 ( .A(n556), .B(n555), .ZN(n683) );
  NAND2_X1 U649 ( .A1(n683), .A2(n557), .ZN(n559) );
  XNOR2_X1 U650 ( .A(KEYINPUT13), .B(G475), .ZN(n558) );
  XNOR2_X1 U651 ( .A(n559), .B(n558), .ZN(n561) );
  INV_X1 U652 ( .A(n561), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n560), .A2(n582), .ZN(n637) );
  NAND2_X1 U654 ( .A1(n583), .A2(n561), .ZN(n728) );
  OR2_X1 U655 ( .A1(n728), .A2(n713), .ZN(n562) );
  XNOR2_X1 U656 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n563) );
  BUF_X1 U657 ( .A(n565), .Z(n711) );
  OR2_X1 U658 ( .A1(n586), .A2(n618), .ZN(n566) );
  OR2_X1 U659 ( .A1(n711), .A2(n566), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n567), .B(KEYINPUT81), .ZN(n568) );
  NAND2_X1 U661 ( .A1(n589), .A2(n568), .ZN(n569) );
  XNOR2_X1 U662 ( .A(n569), .B(KEYINPUT32), .ZN(n775) );
  INV_X1 U663 ( .A(n599), .ZN(n570) );
  AND2_X1 U664 ( .A1(n711), .A2(n347), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n589), .A2(n571), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n572), .B(KEYINPUT65), .ZN(n573) );
  INV_X1 U667 ( .A(n618), .ZN(n714) );
  NAND2_X1 U668 ( .A1(n594), .A2(KEYINPUT44), .ZN(n592) );
  INV_X1 U669 ( .A(KEYINPUT31), .ZN(n576) );
  NOR2_X2 U670 ( .A1(n615), .A2(n710), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n598), .A2(n347), .ZN(n581) );
  AND2_X1 U672 ( .A1(n583), .A2(n582), .ZN(n705) );
  INV_X1 U673 ( .A(n705), .ZN(n666) );
  OR2_X1 U674 ( .A1(n583), .A2(n582), .ZN(n698) );
  AND2_X1 U675 ( .A1(n666), .A2(n698), .ZN(n730) );
  INV_X1 U676 ( .A(n730), .ZN(n630) );
  INV_X1 U677 ( .A(KEYINPUT101), .ZN(n584) );
  XNOR2_X1 U678 ( .A(n585), .B(n584), .ZN(n590) );
  NOR2_X1 U679 ( .A1(n586), .A2(n714), .ZN(n587) );
  AND2_X1 U680 ( .A1(n711), .A2(n587), .ZN(n588) );
  NAND2_X1 U681 ( .A1(n589), .A2(n588), .ZN(n694) );
  AND2_X1 U682 ( .A1(n590), .A2(n694), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U684 ( .A(n593), .B(KEYINPUT89), .ZN(n596) );
  OR2_X1 U685 ( .A1(n594), .A2(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U687 ( .A1(n570), .A2(n725), .ZN(n602) );
  XNOR2_X1 U688 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n600) );
  XNOR2_X1 U689 ( .A(n600), .B(KEYINPUT107), .ZN(n601) );
  XNOR2_X1 U690 ( .A(n602), .B(n601), .ZN(n609) );
  NOR2_X1 U691 ( .A1(G900), .A2(n603), .ZN(n604) );
  NAND2_X1 U692 ( .A1(G953), .A2(n604), .ZN(n605) );
  XNOR2_X1 U693 ( .A(n605), .B(KEYINPUT104), .ZN(n607) );
  AND2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n616) );
  INV_X1 U695 ( .A(n616), .ZN(n608) );
  AND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n633) );
  XOR2_X1 U697 ( .A(KEYINPUT38), .B(n635), .Z(n726) );
  AND2_X1 U698 ( .A1(n633), .A2(n726), .ZN(n610) );
  NAND2_X1 U699 ( .A1(n634), .A2(n610), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n649), .A2(n705), .ZN(n613) );
  XOR2_X1 U701 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n612) );
  NAND2_X1 U702 ( .A1(n726), .A2(n725), .ZN(n729) );
  NOR2_X1 U703 ( .A1(n729), .A2(n728), .ZN(n614) );
  XNOR2_X1 U704 ( .A(KEYINPUT41), .B(n614), .ZN(n739) );
  XNOR2_X1 U705 ( .A(n615), .B(KEYINPUT109), .ZN(n620) );
  NOR2_X1 U706 ( .A1(n739), .A2(n628), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n621), .B(KEYINPUT42), .ZN(n776) );
  NOR2_X2 U708 ( .A1(n673), .A2(n776), .ZN(n622) );
  XNOR2_X1 U709 ( .A(n624), .B(KEYINPUT105), .ZN(n625) );
  XOR2_X1 U710 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n627) );
  NOR2_X1 U711 ( .A1(n632), .A2(KEYINPUT47), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n670), .A2(n631), .ZN(n641) );
  AND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n639) );
  INV_X1 U714 ( .A(n635), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n661) );
  XOR2_X1 U717 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n643) );
  INV_X1 U718 ( .A(n644), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n711), .A2(n725), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT43), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n648), .A2(n635), .ZN(n662) );
  BUF_X1 U723 ( .A(n649), .Z(n650) );
  INV_X1 U724 ( .A(n650), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n651), .A2(n698), .ZN(n663) );
  INV_X1 U726 ( .A(KEYINPUT2), .ZN(n653) );
  INV_X1 U727 ( .A(KEYINPUT64), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n689), .A2(G472), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n767), .A2(G952), .ZN(n659) );
  XOR2_X1 U730 ( .A(G143), .B(KEYINPUT115), .Z(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(G45) );
  XOR2_X1 U732 ( .A(G140), .B(n662), .Z(G42) );
  XOR2_X1 U733 ( .A(G134), .B(n663), .Z(G36) );
  XNOR2_X1 U734 ( .A(G110), .B(KEYINPUT114), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(G12) );
  NOR2_X1 U736 ( .A1(n668), .A2(n666), .ZN(n667) );
  XOR2_X1 U737 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U738 ( .A1(n668), .A2(n698), .ZN(n669) );
  XOR2_X1 U739 ( .A(G116), .B(n669), .Z(G18) );
  XOR2_X1 U740 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(G125), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n670), .B(n672), .ZN(G27) );
  BUF_X1 U743 ( .A(n673), .Z(n674) );
  XOR2_X1 U744 ( .A(n674), .B(G131), .Z(G33) );
  XOR2_X1 U745 ( .A(n675), .B(G122), .Z(G24) );
  NAND2_X1 U746 ( .A1(n689), .A2(G217), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT123), .B(n676), .Z(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U749 ( .A1(n679), .A2(n693), .ZN(G66) );
  NAND2_X1 U750 ( .A1(n689), .A2(G478), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n689), .A2(G475), .ZN(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n689), .A2(G469), .ZN(n688) );
  XNOR2_X1 U754 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT58), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n689), .A2(G210), .ZN(n692) );
  XOR2_X1 U757 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n690) );
  XOR2_X1 U758 ( .A(G101), .B(n694), .Z(n695) );
  XNOR2_X1 U759 ( .A(n695), .B(KEYINPUT113), .ZN(G3) );
  NAND2_X1 U760 ( .A1(n420), .A2(n705), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n697), .B(G104), .ZN(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  INV_X1 U763 ( .A(n698), .ZN(n702) );
  NAND2_X1 U764 ( .A1(n420), .A2(n702), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(G107), .B(n701), .ZN(G9) );
  XOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .Z(n704) );
  NAND2_X1 U768 ( .A1(n702), .A2(n706), .ZN(n703) );
  XNOR2_X1 U769 ( .A(n704), .B(n703), .ZN(G30) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n707), .B(KEYINPUT116), .ZN(n708) );
  XNOR2_X1 U772 ( .A(G146), .B(n708), .ZN(G48) );
  NOR2_X1 U773 ( .A1(n709), .A2(n347), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n712), .B(KEYINPUT50), .ZN(n718) );
  NAND2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U777 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n715) );
  XNOR2_X1 U778 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U780 ( .A(KEYINPUT51), .B(n719), .Z(n720) );
  NOR2_X1 U781 ( .A1(n720), .A2(n570), .ZN(n721) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U783 ( .A1(n723), .A2(n739), .ZN(n735) );
  NOR2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U788 ( .A1(n453), .A2(n733), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(KEYINPUT52), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n742) );
  INV_X1 U792 ( .A(n739), .ZN(n740) );
  AND2_X1 U793 ( .A1(n740), .A2(n724), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n742), .A2(n741), .ZN(n751) );
  NOR2_X1 U795 ( .A1(n757), .A2(KEYINPUT2), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n749) );
  NOR2_X1 U797 ( .A1(n656), .A2(KEYINPUT2), .ZN(n747) );
  INV_X1 U798 ( .A(KEYINPUT86), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U802 ( .A1(n752), .A2(G953), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n753), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U804 ( .A(n754), .B(KEYINPUT125), .ZN(n756) );
  NOR2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n764) );
  NAND2_X1 U806 ( .A1(n757), .A2(n767), .ZN(n762) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n759), .A2(G898), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n760), .B(KEYINPUT124), .ZN(n761) );
  NAND2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U812 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U813 ( .A(n765), .B(n766), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n656), .B(n769), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(n774) );
  XOR2_X1 U816 ( .A(G227), .B(n769), .Z(n770) );
  XNOR2_X1 U817 ( .A(n770), .B(KEYINPUT126), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n774), .A2(n773), .ZN(G72) );
  XNOR2_X1 U821 ( .A(G119), .B(n775), .ZN(G21) );
  XOR2_X1 U822 ( .A(G137), .B(n776), .Z(G39) );
endmodule

