//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n187), .A2(new_n188), .A3(G953), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G122), .ZN(new_n191));
  AOI21_X1  g005(.A(KEYINPUT14), .B1(new_n191), .B2(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(G116), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT92), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G122), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(G122), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n195), .B(new_n197), .C1(new_n198), .C2(KEYINPUT14), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n199), .C1(KEYINPUT14), .C2(new_n197), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n200), .A2(KEYINPUT93), .A3(G107), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT93), .B1(new_n200), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G134), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n198), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n197), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n201), .A2(new_n202), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n212), .B2(new_n197), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n198), .A2(new_n193), .A3(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(KEYINPUT13), .A3(G128), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT91), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT13), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n204), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n204), .A2(new_n222), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT91), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n206), .B(new_n220), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n219), .B1(new_n226), .B2(G134), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n190), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n200), .A2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n200), .A2(KEYINPUT93), .A3(G107), .ZN(new_n232));
  INV_X1    g046(.A(new_n215), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n227), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n189), .ZN(new_n236));
  AOI21_X1  g050(.A(G902), .B1(new_n228), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G478), .ZN(new_n239));
  OR3_X1    g053(.A1(new_n237), .A2(KEYINPUT94), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT94), .B1(new_n237), .B2(new_n239), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n216), .A2(new_n227), .A3(new_n190), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n189), .B1(new_n234), .B2(new_n235), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n239), .B(KEYINPUT95), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n242), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n237), .A2(KEYINPUT96), .A3(new_n247), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n240), .A2(new_n241), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n254), .B2(KEYINPUT88), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(KEYINPUT88), .B2(new_n254), .ZN(new_n256));
  XNOR2_X1  g070(.A(G113), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(G104), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n260));
  INV_X1    g074(.A(G140), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G140), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT19), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G125), .B(G140), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT19), .ZN(new_n269));
  AOI21_X1  g083(.A(G146), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n263), .A2(KEYINPUT16), .A3(G140), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT16), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n272), .A2(new_n273), .A3(G146), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n260), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G237), .A2(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G214), .ZN(new_n277));
  OR2_X1    g091(.A1(KEYINPUT84), .A2(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT84), .A2(G143), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n277), .A2(new_n279), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(G214), .A3(new_n276), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n279), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n271), .B1(new_n268), .B2(KEYINPUT16), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G146), .ZN(new_n290));
  INV_X1    g104(.A(G146), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT19), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT19), .B1(new_n262), .B2(new_n264), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT85), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n275), .A2(new_n288), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n265), .A2(G146), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n268), .A2(new_n291), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n286), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT18), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(new_n285), .ZN(new_n302));
  OAI221_X1 g116(.A(new_n299), .B1(new_n300), .B2(new_n302), .C1(new_n282), .C2(new_n301), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n296), .A2(new_n303), .A3(KEYINPUT86), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n259), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n282), .A2(new_n309), .A3(new_n287), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT87), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n289), .A2(G146), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(new_n274), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT87), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n282), .A2(new_n287), .A3(new_n314), .A4(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(KEYINPUT17), .A3(G131), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n313), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n303), .A3(new_n259), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n256), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n253), .B1(new_n308), .B2(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT20), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT89), .B(new_n256), .C1(new_n308), .C2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n303), .ZN(new_n327));
  INV_X1    g141(.A(new_n259), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n243), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g145(.A(G475), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(G234), .A2(G237), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(G952), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT21), .B(G898), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(G902), .A3(G953), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n251), .A2(new_n326), .A3(new_n332), .A4(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G214), .B1(G237), .B2(G902), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT2), .B(G113), .Z(new_n342));
  XNOR2_X1  g156(.A(G116), .B(G119), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n196), .A2(KEYINPUT5), .A3(G119), .ZN(new_n346));
  INV_X1    g160(.A(G113), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n213), .A2(G104), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n258), .A2(G107), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n258), .B2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(KEYINPUT3), .C1(new_n258), .C2(G107), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n353), .B1(new_n359), .B2(new_n350), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n349), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n213), .A2(G104), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n258), .A2(G107), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n357), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(new_n358), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n365), .B(new_n350), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n358), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n370), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT78), .B1(new_n370), .B2(new_n365), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n373), .B2(G101), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n365), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n359), .A2(KEYINPUT78), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n342), .A2(new_n343), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n344), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n361), .B1(new_n374), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G122), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n361), .B(new_n386), .C1(new_n374), .C2(new_n384), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n291), .A2(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n203), .A2(G146), .ZN(new_n394));
  AOI21_X1  g208(.A(G128), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n203), .A2(KEYINPUT1), .A3(G146), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT66), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n399));
  XNOR2_X1  g213(.A(G143), .B(G146), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n399), .B(new_n396), .C1(new_n400), .C2(G128), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n393), .A2(new_n394), .A3(new_n402), .A4(G128), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n263), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT64), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G128), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n393), .A2(new_n394), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n205), .A2(KEYINPUT0), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT0), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n413), .A3(KEYINPUT64), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n400), .A2(new_n416), .A3(KEYINPUT0), .A4(G128), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n400), .A2(KEYINPUT0), .A3(G128), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT65), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n415), .A2(G125), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n405), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n334), .A2(G224), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT82), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n421), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n390), .A2(new_n392), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n405), .A2(new_n420), .A3(KEYINPUT83), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n386), .B(KEYINPUT8), .ZN(new_n430));
  INV_X1    g244(.A(new_n361), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n349), .A2(new_n360), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n434));
  INV_X1    g248(.A(new_n428), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n421), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n421), .A2(new_n435), .ZN(new_n437));
  AND4_X1   g251(.A1(new_n429), .A2(new_n433), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n438), .B2(new_n389), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n426), .A2(new_n427), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n427), .B1(new_n426), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n341), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n340), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n209), .B2(G137), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n209), .A2(G137), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n448), .A3(new_n285), .A4(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n415), .A2(new_n452), .A3(new_n417), .A4(new_n419), .ZN(new_n453));
  INV_X1    g267(.A(new_n446), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n209), .A2(G137), .ZN(new_n455));
  OAI21_X1  g269(.A(G131), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n451), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n404), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n459), .A3(new_n382), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n382), .B1(new_n453), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT28), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n276), .A2(G210), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT27), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT26), .B(G101), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND4_X1   g286(.A1(new_n452), .A2(new_n415), .A3(new_n417), .A4(new_n419), .ZN(new_n473));
  AND4_X1   g287(.A1(new_n402), .A2(new_n393), .A3(new_n394), .A4(G128), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n396), .B1(new_n400), .B2(G128), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(KEYINPUT66), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n457), .B1(new_n476), .B2(new_n401), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT30), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n453), .A2(new_n459), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n461), .B1(new_n481), .B2(new_n383), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n467), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n472), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n243), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  OAI21_X1  g300(.A(G472), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT67), .B(KEYINPUT31), .Z(new_n489));
  NAND4_X1  g303(.A1(new_n482), .A2(KEYINPUT68), .A3(new_n467), .A4(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n453), .A2(new_n459), .A3(new_n479), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n453), .B2(new_n459), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n383), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n493), .A2(new_n460), .A3(new_n467), .A4(new_n489), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n460), .A3(new_n467), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n467), .B1(new_n463), .B2(new_n469), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(KEYINPUT31), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n488), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n502), .ZN(new_n504));
  AOI211_X1 g318(.A(KEYINPUT32), .B(new_n504), .C1(new_n497), .C2(new_n500), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n487), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n476), .B2(new_n401), .ZN(new_n510));
  INV_X1    g324(.A(new_n353), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n403), .B(new_n396), .C1(G128), .C2(new_n400), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n368), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n510), .A2(new_n360), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n415), .A2(new_n417), .A3(new_n419), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n380), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n374), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n452), .ZN(new_n518));
  INV_X1    g332(.A(new_n452), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n514), .B(new_n519), .C1(new_n374), .C2(new_n516), .ZN(new_n520));
  XNOR2_X1  g334(.A(G110), .B(G140), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT76), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n334), .A2(G227), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n513), .B1(new_n360), .B2(new_n404), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n452), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(KEYINPUT12), .A3(new_n452), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n520), .ZN(new_n532));
  INV_X1    g346(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT79), .B1(new_n531), .B2(new_n520), .ZN(new_n535));
  OAI211_X1 g349(.A(G469), .B(new_n525), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G469), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n243), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n520), .A2(new_n524), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT80), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n520), .A2(new_n543), .A3(new_n524), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n544), .A3(new_n531), .ZN(new_n545));
  INV_X1    g359(.A(new_n520), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n371), .A2(new_n372), .A3(new_n350), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n515), .B(new_n380), .C1(new_n547), .C2(new_n369), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n519), .B1(new_n548), .B2(new_n514), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n533), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n518), .A2(new_n520), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT81), .A3(new_n533), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n537), .A3(new_n243), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n508), .B1(new_n540), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT70), .B1(new_n205), .B2(G119), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  INV_X1    g373(.A(G119), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(G128), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n558), .B(new_n561), .C1(new_n560), .C2(G128), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n560), .B2(G128), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n560), .A2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(G110), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n290), .B(new_n298), .C1(new_n564), .C2(new_n570), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n312), .A2(new_n274), .B1(new_n563), .B2(new_n562), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(KEYINPUT71), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n569), .A2(KEYINPUT71), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n571), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT73), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n571), .B(new_n579), .C1(new_n572), .C2(new_n576), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT72), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT22), .B(G137), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n577), .A2(KEYINPUT73), .A3(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(G217), .A2(G902), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n188), .B2(G234), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(KEYINPUT69), .Z(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n585), .B2(new_n586), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT25), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT74), .B(KEYINPUT25), .Z(new_n597));
  AOI211_X1 g411(.A(G902), .B(new_n597), .C1(new_n585), .C2(new_n586), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n592), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT75), .B(new_n592), .C1(new_n596), .C2(new_n598), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n443), .A2(new_n506), .A3(new_n557), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI21_X1  g419(.A(new_n383), .B1(new_n473), .B2(new_n477), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n468), .B1(new_n606), .B2(new_n460), .ZN(new_n607));
  INV_X1    g421(.A(new_n469), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n484), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT31), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n496), .A2(new_n490), .B1(new_n611), .B2(new_n498), .ZN(new_n612));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT97), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n612), .A2(G902), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n614), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n501), .B2(new_n243), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n557), .A2(new_n618), .A3(new_n603), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n426), .A2(new_n439), .ZN(new_n620));
  INV_X1    g434(.A(new_n427), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n426), .A2(new_n439), .A3(new_n427), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n341), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n441), .B2(KEYINPUT98), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n296), .A2(new_n303), .A3(KEYINPUT86), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT86), .B1(new_n296), .B2(new_n303), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n328), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n254), .B1(new_n631), .B2(new_n318), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n325), .B1(new_n252), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n318), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT89), .B1(new_n634), .B2(new_n256), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n332), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n237), .B2(G478), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  INV_X1    g452(.A(G478), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n246), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n244), .B2(new_n245), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n228), .A2(new_n644), .A3(new_n236), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n639), .A2(G902), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n647), .ZN(new_n649));
  AOI211_X1 g463(.A(KEYINPUT99), .B(new_n649), .C1(new_n643), .C2(new_n645), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n641), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n636), .A2(new_n651), .A3(new_n339), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n619), .A2(new_n628), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT34), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  OR3_X1    g469(.A1(new_n632), .A2(KEYINPUT101), .A3(new_n252), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n332), .ZN(new_n657));
  INV_X1    g471(.A(new_n251), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n339), .B(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n632), .A2(new_n252), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n324), .A2(new_n660), .A3(KEYINPUT101), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  OR3_X1    g476(.A1(new_n662), .A2(new_n628), .A3(KEYINPUT103), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n662), .B2(new_n628), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n619), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT35), .B(G107), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n584), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n577), .B(new_n669), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n591), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n596), .B2(new_n598), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n443), .A2(new_n618), .A3(new_n557), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR3_X1   g489(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n620), .A2(KEYINPUT98), .A3(new_n621), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n341), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n506), .A3(new_n557), .A4(new_n672), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n338), .A2(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n335), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n657), .A2(new_n658), .A3(new_n661), .A4(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n205), .ZN(G30));
  NOR2_X1   g499(.A1(new_n440), .A2(new_n441), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT38), .Z(new_n687));
  AND4_X1   g501(.A1(new_n341), .A2(new_n687), .A3(new_n636), .A4(new_n658), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n540), .A2(new_n556), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n507), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n682), .B(KEYINPUT39), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT40), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT32), .B1(new_n612), .B2(new_n504), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n501), .A2(new_n488), .A3(new_n502), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n482), .A2(new_n484), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n461), .A2(new_n462), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n698), .B2(new_n484), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n672), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OR3_X1    g519(.A1(new_n690), .A2(KEYINPUT40), .A3(new_n692), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n688), .A2(new_n693), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND3_X1  g522(.A1(new_n636), .A2(new_n651), .A3(new_n682), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n636), .A2(new_n651), .A3(KEYINPUT104), .A4(new_n682), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n680), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n291), .ZN(G48));
  NAND2_X1  g529(.A1(new_n556), .A2(new_n507), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT81), .B1(new_n553), .B2(new_n533), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n551), .B(new_n524), .C1(new_n518), .C2(new_n520), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(G902), .B1(new_n719), .B2(new_n545), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT105), .B1(new_n720), .B2(new_n537), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n555), .A2(new_n243), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(G469), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n716), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n601), .A2(new_n602), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n696), .B2(new_n487), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n628), .A2(new_n652), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n721), .A2(new_n724), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n508), .B1(new_n720), .B2(new_n537), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n663), .B2(new_n664), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n196), .ZN(G18));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n723), .B1(new_n722), .B2(G469), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT105), .B(new_n537), .C1(new_n555), .C2(new_n243), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n737), .B1(new_n740), .B2(new_n628), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n679), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n506), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n340), .A3(new_n703), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n560), .ZN(G21));
  NAND2_X1  g561(.A1(new_n658), .A2(new_n636), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n628), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n725), .A2(new_n659), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT107), .B1(new_n612), .B2(new_n504), .ZN(new_n752));
  OAI21_X1  g566(.A(G472), .B1(new_n612), .B2(G902), .ZN(new_n753));
  INV_X1    g567(.A(new_n599), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n501), .A2(new_n755), .A3(new_n502), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT108), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n191), .ZN(G24));
  AND4_X1   g574(.A1(new_n672), .A2(new_n752), .A3(new_n753), .A4(new_n756), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n711), .A3(new_n712), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n741), .B2(new_n742), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n263), .ZN(G27));
  AND2_X1   g578(.A1(new_n711), .A2(new_n712), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n440), .A2(new_n441), .A3(new_n626), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n557), .A2(KEYINPUT42), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n599), .B1(new_n696), .B2(new_n487), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n506), .A2(new_n557), .A3(new_n603), .A4(new_n766), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n713), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n683), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n209), .ZN(G36));
  OAI21_X1  g590(.A(new_n525), .B1(new_n534), .B2(new_n535), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n537), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n525), .C1(new_n534), .C2(new_n535), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n538), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n556), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n507), .B(new_n691), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n618), .A2(new_n703), .ZN(new_n787));
  INV_X1    g601(.A(new_n636), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n651), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n651), .B1(KEYINPUT111), .B2(KEYINPUT43), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n788), .C1(KEYINPUT111), .C2(new_n651), .ZN(new_n792));
  OR2_X1    g606(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n787), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n766), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n784), .A2(new_n785), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n786), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NOR2_X1   g615(.A1(new_n797), .A2(new_n603), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n765), .A2(new_n744), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n507), .B1(new_n782), .B2(new_n783), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT112), .B(new_n507), .C1(new_n782), .C2(new_n783), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n804), .B(KEYINPUT47), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n804), .A2(KEYINPUT47), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n805), .B2(new_n806), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n804), .A2(KEYINPUT47), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n808), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n803), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n261), .ZN(G42));
  NAND3_X1  g630(.A1(new_n732), .A2(new_n508), .A3(new_n556), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n335), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n819), .A2(new_n790), .A3(new_n792), .A4(new_n793), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n341), .A2(new_n820), .A3(new_n686), .A4(new_n758), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n818), .A2(new_n824), .A3(new_n821), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n687), .A2(new_n341), .A3(new_n740), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n820), .A3(new_n758), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n827), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n740), .A2(new_n797), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n820), .A2(new_n761), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n702), .A2(new_n726), .A3(new_n335), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n636), .A2(new_n651), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n830), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n823), .A2(new_n825), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n820), .A2(new_n768), .A3(new_n831), .ZN(new_n841));
  XNOR2_X1  g655(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n844));
  INV_X1    g658(.A(G952), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n636), .A2(new_n651), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n845), .B(G953), .C1(new_n834), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n743), .A2(new_n758), .A3(new_n820), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n844), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n836), .A2(new_n832), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n827), .A2(KEYINPUT118), .A3(new_n828), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n827), .B1(KEYINPUT118), .B2(new_n828), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n851), .B(KEYINPUT51), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n850), .B1(new_n855), .B2(new_n822), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n775), .B1(new_n769), .B2(new_n772), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n557), .A2(new_n766), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n762), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n860), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n765), .A2(new_n862), .A3(KEYINPUT116), .A4(new_n761), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n744), .A2(new_n703), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n251), .A2(new_n657), .A3(new_n661), .A4(new_n682), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n858), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n341), .B(new_n659), .C1(new_n440), .C2(new_n441), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n636), .A3(new_n251), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n603), .A3(new_n618), .A4(new_n557), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n729), .A2(new_n673), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n735), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n743), .A2(new_n745), .B1(new_n751), .B2(new_n758), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n846), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n603), .A3(new_n557), .A4(new_n618), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n876), .A2(new_n604), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n876), .B2(new_n604), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n868), .A2(new_n873), .A3(new_n874), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n762), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n740), .A2(new_n737), .A3(new_n628), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT106), .B1(new_n725), .B2(new_n679), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n680), .B1(new_n683), .B2(new_n713), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n788), .A2(new_n251), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n679), .A2(new_n888), .A3(new_n557), .A4(new_n682), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n704), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n743), .B2(new_n882), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n857), .B1(new_n881), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n895), .B1(new_n894), .B2(new_n891), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n763), .A2(new_n886), .A3(KEYINPUT52), .A4(new_n890), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n874), .A2(new_n873), .A3(new_n880), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n858), .A2(new_n864), .A3(new_n867), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT53), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n898), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n898), .B2(new_n905), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n840), .B(new_n856), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n845), .A2(new_n334), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n754), .A2(new_n507), .A3(new_n341), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n732), .A2(new_n556), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n789), .B(new_n911), .C1(new_n912), .C2(KEYINPUT49), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT114), .Z(new_n914));
  NOR2_X1   g728(.A1(new_n687), .A2(new_n702), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n915), .C1(KEYINPUT49), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n916), .ZN(G75));
  NOR3_X1   g731(.A1(new_n881), .A2(new_n897), .A3(new_n857), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n901), .B2(new_n904), .ZN(new_n919));
  OAI211_X1 g733(.A(G210), .B(G902), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n390), .A2(new_n392), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n425), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n920), .B2(new_n921), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n334), .A2(G952), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G51));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n918), .B2(new_n919), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n898), .A2(new_n905), .A3(KEYINPUT54), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n538), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n555), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n243), .B1(new_n898), .B2(new_n905), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n780), .A3(new_n779), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n928), .B1(new_n936), .B2(new_n938), .ZN(G54));
  AND2_X1   g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n631), .A3(new_n318), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n634), .A3(new_n940), .ZN(new_n943));
  INV_X1    g757(.A(new_n928), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G60));
  NOR2_X1   g759(.A1(new_n906), .A2(new_n907), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n646), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n931), .A2(new_n646), .A3(new_n932), .A4(new_n948), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G63));
  INV_X1    g766(.A(new_n587), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n918), .A2(new_n919), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n588), .B(KEYINPUT60), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n898), .B2(new_n905), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n928), .B1(new_n957), .B2(new_n670), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n957), .B2(new_n670), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n956), .B(new_n958), .C1(new_n960), .C2(KEYINPUT61), .ZN(new_n961));
  INV_X1    g775(.A(new_n955), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n670), .B(new_n962), .C1(new_n918), .C2(new_n919), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n963), .B(new_n944), .C1(new_n587), .C2(new_n957), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT61), .B1(new_n963), .B2(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n966), .ZN(G66));
  AOI21_X1  g781(.A(new_n334), .B1(new_n337), .B2(G224), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n902), .B2(new_n334), .ZN(new_n969));
  INV_X1    g783(.A(G898), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n922), .B1(new_n970), .B2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n969), .B(new_n971), .ZN(G69));
  OAI21_X1  g786(.A(new_n846), .B1(new_n636), .B2(new_n251), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(new_n727), .A3(new_n691), .A4(new_n862), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n800), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n803), .ZN(new_n977));
  INV_X1    g791(.A(new_n814), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n813), .B1(new_n812), .B2(new_n808), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n707), .A2(new_n894), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n707), .A2(new_n894), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n976), .A2(new_n980), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n334), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n292), .A2(new_n293), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n481), .B(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n786), .A2(new_n749), .A3(new_n768), .A4(new_n799), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n800), .A2(new_n989), .A3(new_n858), .A4(new_n894), .ZN(new_n990));
  OR3_X1    g804(.A1(new_n990), .A2(new_n815), .A3(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(G900), .B2(G953), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n986), .A2(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n334), .B1(G227), .B2(G900), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n993), .B(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(new_n482), .A2(new_n484), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT127), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n990), .A2(new_n815), .A3(new_n902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n613), .A2(new_n243), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n697), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1003), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n998), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n944), .B(new_n1004), .C1(new_n954), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n985), .B2(new_n902), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n697), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(G57));
endmodule


