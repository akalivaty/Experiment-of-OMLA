//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  NOR3_X1   g000(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT27), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G183gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n213), .C1(new_n214), .C2(new_n211), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n212), .A2(KEYINPUT67), .A3(KEYINPUT68), .A4(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT28), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n214), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n219));
  OAI221_X1 g018(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(new_n208), .B2(new_n209), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n225), .B(KEYINPUT64), .ZN(new_n235));
  NOR4_X1   g034(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT25), .A4(new_n232), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n234), .A2(KEYINPUT25), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n239), .B2(G134gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT71), .B(new_n240), .C1(new_n241), .C2(KEYINPUT70), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT70), .A2(KEYINPUT71), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(new_n239), .A3(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G113gat), .B(G120gat), .Z(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(KEYINPUT72), .A3(new_n244), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n253));
  NAND2_X1  g052(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n248), .A2(new_n241), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n238), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n256), .A2(new_n220), .A3(new_n237), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n257), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT34), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n262), .A3(new_n260), .ZN(new_n266));
  INV_X1    g065(.A(new_n261), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT32), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(KEYINPUT33), .ZN(new_n269));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G71gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G99gat), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n268), .B(new_n277), .C1(new_n266), .C2(new_n267), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n265), .A2(new_n273), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n269), .A2(new_n272), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n264), .B1(new_n281), .B2(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(KEYINPUT36), .A3(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT76), .B(G218gat), .Z(new_n288));
  INV_X1    g087(.A(G211gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G211gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n289), .A3(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G141gat), .B(G148gat), .Z(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT2), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT3), .B1(new_n297), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(G22gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G78gat), .B(G106gat), .Z(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT31), .ZN(new_n319));
  INV_X1    g118(.A(G50gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT81), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n310), .B(new_n315), .C1(new_n311), .C2(new_n305), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n322), .A2(KEYINPUT81), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(KEYINPUT82), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n317), .A2(new_n327), .A3(new_n323), .A4(new_n324), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n329), .A2(KEYINPUT83), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT83), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n256), .A2(new_n340), .A3(new_n305), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n252), .A2(new_n305), .A3(new_n255), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n252), .A2(new_n255), .B1(new_n306), .B2(KEYINPUT3), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n341), .A2(new_n343), .B1(new_n307), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n257), .A2(new_n306), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n339), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT5), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n338), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n339), .ZN(new_n355));
  INV_X1    g154(.A(new_n338), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(new_n348), .B2(new_n342), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n345), .B2(new_n346), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n355), .B(new_n356), .C1(new_n358), .C2(new_n339), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n352), .A2(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  INV_X1    g164(.A(G64gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT77), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n238), .B2(new_n308), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(KEYINPUT78), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(new_n220), .B2(new_n237), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n297), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n238), .A2(new_n371), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n220), .B2(new_n237), .ZN(new_n377));
  INV_X1    g176(.A(new_n373), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n298), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n380), .A2(KEYINPUT30), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n369), .B(KEYINPUT79), .Z(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(KEYINPUT30), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n364), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n285), .A2(new_n286), .B1(new_n333), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n329), .A2(new_n330), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n379), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT37), .A3(new_n379), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n369), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n380), .B1(new_n393), .B2(KEYINPUT38), .ZN(new_n394));
  OR3_X1    g193(.A1(new_n372), .A2(new_n374), .A3(new_n297), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n377), .A2(new_n378), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n238), .B2(new_n371), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(KEYINPUT37), .C1(new_n397), .C2(new_n298), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT38), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n382), .A4(new_n391), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n394), .A2(new_n363), .A3(new_n361), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n345), .A2(KEYINPUT39), .A3(new_n346), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n356), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n341), .A2(new_n343), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n344), .A2(new_n307), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n350), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT84), .B(new_n338), .C1(new_n408), .C2(KEYINPUT39), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n408), .B(KEYINPUT39), .C1(new_n350), .C2(new_n349), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT40), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(KEYINPUT40), .A3(new_n411), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT40), .B1(new_n410), .B2(new_n411), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n359), .B1(new_n419), .B2(new_n413), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n388), .B(new_n401), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n387), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n280), .A2(new_n388), .A3(new_n282), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n416), .B1(new_n363), .B2(new_n361), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT35), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT35), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n386), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G15gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n314), .ZN(new_n432));
  NAND2_X1  g231(.A1(G15gat), .A2(G22gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT90), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT16), .B1(new_n432), .B2(new_n433), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n436), .A2(G1gat), .A3(G8gat), .ZN(new_n437));
  INV_X1    g236(.A(G8gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT16), .ZN(new_n439));
  AND2_X1   g238(.A1(G15gat), .A2(G22gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(G15gat), .A2(G22gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G1gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n435), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(G8gat), .B1(new_n436), .B2(G1gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n435), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n443), .A3(new_n438), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n320), .A2(G43gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT15), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n320), .A2(G43gat), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G29gat), .ZN(new_n457));
  INV_X1    g256(.A(G36gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT87), .B1(new_n320), .B2(G43gat), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461));
  INV_X1    g260(.A(G43gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(G50gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n463), .A3(new_n451), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n464), .B2(new_n453), .ZN(new_n465));
  OAI22_X1  g264(.A1(KEYINPUT86), .A2(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND4_X1   g268(.A1(KEYINPUT86), .A2(new_n457), .A3(new_n458), .A4(KEYINPUT14), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(new_n468), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT88), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n456), .B(new_n465), .C1(new_n472), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n475), .B(new_n476), .C1(new_n457), .C2(new_n458), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n455), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT17), .B1(new_n481), .B2(KEYINPUT89), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n484));
  AOI211_X1 g283(.A(new_n483), .B(new_n484), .C1(new_n478), .C2(new_n480), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n450), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n471), .B1(new_n469), .B2(new_n470), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT88), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n455), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n489), .A2(new_n465), .B1(new_n479), .B2(new_n455), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT91), .B1(new_n490), .B2(new_n450), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n437), .A2(new_n444), .A3(new_n435), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n481), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n486), .A2(KEYINPUT18), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n490), .A2(new_n450), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n490), .A2(new_n450), .A3(KEYINPUT91), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n494), .B2(new_n481), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n498), .B(KEYINPUT13), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT93), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G197gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT11), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(new_n230), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n499), .A2(new_n506), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n486), .A2(new_n497), .A3(new_n498), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT92), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n486), .A2(new_n519), .A3(new_n497), .A4(new_n498), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n514), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n514), .B1(new_n515), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(G85gat), .A3(G92gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n525), .A2(new_n528), .A3(G85gat), .A4(G92gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT101), .B(G85gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n368), .ZN(new_n532));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT8), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n533), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n530), .A2(new_n532), .A3(new_n538), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n482), .B2(new_n485), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n481), .A2(new_n539), .A3(new_n537), .ZN(new_n542));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT98), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT41), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G190gat), .B(G218gat), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n541), .A2(new_n548), .A3(new_n542), .A4(new_n546), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT99), .B(G134gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G162gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n544), .A2(new_n545), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(KEYINPUT102), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n559), .A2(new_n555), .B1(new_n550), .B2(new_n551), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n565), .B2(KEYINPUT94), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n562), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G64gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n366), .A2(G57gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n570), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(KEYINPUT9), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  NOR2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT95), .A4(new_n566), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n570), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT97), .B1(new_n583), .B2(new_n586), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n595));
  INV_X1    g394(.A(new_n586), .ZN(new_n596));
  AOI211_X1 g395(.A(new_n595), .B(new_n596), .C1(new_n572), .C2(new_n582), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT21), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n598), .A2(new_n600), .A3(new_n450), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(new_n598), .B2(new_n450), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n593), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT20), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n595), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n583), .A2(KEYINPUT97), .A3(new_n586), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n588), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n599), .B1(new_n609), .B2(new_n494), .ZN(new_n610));
  INV_X1    g409(.A(new_n593), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n600), .A3(new_n450), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n603), .A2(new_n606), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n606), .B1(new_n603), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n592), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n603), .A2(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n605), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n613), .A3(new_n606), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n591), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n561), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n561), .A2(new_n616), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n587), .A2(new_n540), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n583), .A2(new_n537), .A3(new_n539), .A4(new_n586), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n537), .A2(KEYINPUT10), .A3(new_n539), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n594), .B2(new_n597), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n626), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n629), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n626), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT104), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n231), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(G204gat), .Z(new_n640));
  OR2_X1    g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n630), .A2(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n625), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n635), .A2(new_n626), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n640), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n622), .A2(new_n624), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT105), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n622), .A2(new_n650), .A3(new_n624), .A4(new_n647), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n524), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n430), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n364), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n443), .ZN(G1324gat));
  AOI211_X1 g454(.A(new_n385), .B(new_n653), .C1(KEYINPUT16), .C2(G8gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n657));
  OAI21_X1  g456(.A(G8gat), .B1(new_n653), .B2(new_n385), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  MUX2_X1   g458(.A(new_n657), .B(new_n659), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g459(.A1(new_n285), .A2(new_n286), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n653), .A2(new_n431), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n431), .B1(new_n653), .B2(new_n283), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(G1326gat));
  INV_X1    g466(.A(new_n333), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  AOI21_X1  g470(.A(new_n561), .B1(new_n422), .B2(new_n429), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT44), .B(new_n561), .C1(new_n422), .C2(new_n429), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n616), .A2(new_n620), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n524), .A3(new_n646), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n364), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n672), .A2(new_n679), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n364), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n457), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT107), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(KEYINPUT45), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(KEYINPUT45), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n681), .B1(new_n687), .B2(new_n688), .ZN(G1328gat));
  OAI21_X1  g488(.A(G36gat), .B1(new_n680), .B2(new_n385), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n682), .A2(G36gat), .A3(new_n385), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT46), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(new_n283), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n683), .A2(new_n462), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n662), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n462), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT47), .B(new_n695), .C1(new_n696), .C2(new_n462), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  OAI21_X1  g500(.A(KEYINPUT108), .B1(new_n680), .B2(new_n388), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  INV_X1    g502(.A(new_n388), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n676), .A2(new_n703), .A3(new_n704), .A4(new_n679), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(G50gat), .A3(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n682), .A2(G50gat), .A3(new_n668), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(KEYINPUT48), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n680), .A2(new_n668), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n710), .B2(new_n320), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n622), .A2(new_n624), .A3(new_n646), .A4(new_n524), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n430), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n364), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n573), .ZN(G1332gat));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n385), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT49), .B(G64gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(G1333gat));
  NOR3_X1   g523(.A1(new_n717), .A2(new_n563), .A3(new_n662), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT110), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n563), .B1(new_n717), .B2(new_n283), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g528(.A1(new_n717), .A2(new_n668), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n564), .ZN(G1335gat));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n559), .A2(new_n555), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n550), .A2(new_n551), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n556), .ZN(new_n736));
  INV_X1    g535(.A(new_n524), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n678), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n732), .A2(new_n430), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n732), .B1(new_n672), .B2(new_n738), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n647), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n684), .A3(new_n531), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n737), .A2(new_n678), .A3(new_n647), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n674), .B2(new_n675), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(KEYINPUT111), .B(new_n746), .C1(new_n674), .C2(new_n675), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n364), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n751), .B2(new_n531), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n430), .A2(new_n736), .A3(new_n738), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT112), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n739), .B2(new_n741), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n416), .A2(new_n368), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n647), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(KEYINPUT112), .A3(new_n732), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n755), .A2(KEYINPUT113), .A3(new_n757), .A4(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n749), .A2(new_n750), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n368), .B1(new_n764), .B2(new_n416), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n747), .B2(new_n385), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(new_n744), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n756), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1337gat));
  AOI21_X1  g570(.A(G99gat), .B1(new_n744), .B2(new_n694), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n662), .B1(new_n749), .B2(new_n750), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(G99gat), .B2(new_n773), .ZN(G1338gat));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n676), .A2(new_n775), .A3(new_n704), .A4(new_n746), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT115), .B1(new_n747), .B2(new_n388), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(G106gat), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n388), .A2(G106gat), .A3(new_n647), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT114), .Z(new_n781));
  OAI211_X1 g580(.A(new_n778), .B(new_n779), .C1(new_n743), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n755), .A2(new_n758), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n781), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n333), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(G106gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n786), .B2(new_n779), .ZN(G1339gat));
  NAND3_X1  g586(.A1(new_n630), .A2(new_n633), .A3(new_n626), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n643), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n640), .B1(new_n634), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT55), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n645), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(new_n789), .B2(new_n791), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n789), .C2(new_n791), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n736), .B(new_n793), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n486), .A2(new_n497), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(G229gat), .A3(G233gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n497), .A2(new_n500), .A3(new_n504), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n511), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n513), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n521), .A2(new_n805), .A3(new_n515), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n645), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n791), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n795), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n521), .A2(new_n515), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n803), .B1(new_n817), .B2(new_n805), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n736), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n646), .A3(new_n806), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n524), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n808), .A2(new_n819), .B1(new_n822), .B2(new_n561), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n823), .A2(new_n678), .B1(new_n648), .B2(new_n737), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n364), .A3(new_n416), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n668), .A3(new_n694), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n524), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n424), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n524), .A2(G113gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n827), .B2(new_n647), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n647), .A2(G120gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n829), .B2(new_n833), .ZN(G1341gat));
  NOR3_X1   g633(.A1(new_n827), .A2(new_n239), .A3(new_n677), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n829), .A2(new_n677), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT118), .Z(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n239), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n829), .A2(G134gat), .A3(new_n561), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT56), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n827), .B2(new_n561), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n808), .A2(new_n819), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n822), .A2(new_n561), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n678), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n648), .A2(new_n737), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n704), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n524), .A2(new_n809), .A3(new_n794), .ZN(new_n851));
  INV_X1    g650(.A(new_n820), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n561), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n843), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n846), .B1(new_n854), .B2(new_n677), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n668), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n661), .A2(new_n364), .A3(new_n416), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n524), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n848), .A2(new_n857), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n860), .A2(G141gat), .A3(new_n524), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(G1344gat));
  INV_X1    g663(.A(new_n860), .ZN(new_n865));
  INV_X1    g664(.A(G148gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n646), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n858), .B2(new_n647), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n866), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n668), .A2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n649), .A2(new_n651), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n524), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n815), .A2(new_n736), .A3(new_n818), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n853), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n677), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n872), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n849), .B1(new_n824), .B2(new_n704), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n646), .A3(new_n857), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n868), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n867), .B1(new_n870), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(new_n300), .B1(new_n860), .B2(new_n677), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n678), .A2(G155gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n858), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT120), .Z(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n858), .B2(new_n561), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n301), .A3(new_n736), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n825), .A2(new_n684), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n424), .A2(KEYINPUT121), .A3(new_n416), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT121), .B1(new_n424), .B2(new_n416), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n230), .A3(new_n737), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n891), .A2(new_n416), .A3(new_n668), .A4(new_n694), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n524), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1348gat));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n231), .A3(new_n646), .ZN(new_n900));
  OAI21_X1  g699(.A(G176gat), .B1(new_n897), .B2(new_n647), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT122), .Z(G1349gat));
  NAND3_X1  g702(.A1(new_n895), .A2(new_n214), .A3(new_n678), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n897), .B2(new_n677), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n897), .B2(new_n561), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT61), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n209), .A3(new_n736), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n661), .A2(new_n684), .A3(new_n385), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n848), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G197gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n737), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n878), .B2(new_n879), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n737), .B1(new_n649), .B2(new_n651), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n678), .B1(new_n853), .B2(new_n875), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n871), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n913), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n737), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n917), .B1(new_n927), .B2(new_n916), .ZN(G1352gat));
  AND3_X1   g727(.A1(new_n919), .A2(new_n923), .A3(new_n922), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n919), .B2(new_n922), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n646), .B(new_n913), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  XOR2_X1   g731(.A(KEYINPUT125), .B(G204gat), .Z(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n925), .A2(new_n934), .A3(new_n646), .A4(new_n913), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n914), .A2(new_n647), .A3(new_n933), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n936), .A2(KEYINPUT127), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n880), .A2(new_n678), .A3(new_n913), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G211gat), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  NAND3_X1  g745(.A1(new_n915), .A2(new_n289), .A3(new_n678), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n915), .B2(new_n736), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n561), .A2(new_n288), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n926), .B2(new_n950), .ZN(G1355gat));
endmodule


