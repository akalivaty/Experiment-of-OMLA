//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT84), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n216), .A3(new_n218), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(KEYINPUT85), .A2(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT85), .A2(KEYINPUT17), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n223), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT85), .A3(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n231), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(G8gat), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n228), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n210), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n235), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n240), .B(KEYINPUT13), .Z(new_n245));
  AOI22_X1  g044(.A1(new_n242), .A2(KEYINPUT18), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n210), .B(new_n247), .C1(new_n239), .C2(new_n241), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n209), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n236), .A2(new_n240), .A3(new_n238), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT18), .B1(new_n250), .B2(KEYINPUT86), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n245), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(new_n209), .A3(new_n248), .A4(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G183gat), .B(G211gat), .ZN(new_n256));
  INV_X1    g055(.A(G155gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT92), .B(G127gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G231gat), .A2(G233gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G64gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G57gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT89), .B(G57gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(new_n266), .ZN(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G78gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT90), .Z(new_n272));
  XOR2_X1   g071(.A(G57gat), .B(G64gat), .Z(new_n273));
  AOI21_X1  g072(.A(new_n270), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT20), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n235), .B1(new_n277), .B2(new_n278), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n280), .B2(new_n282), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n262), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n282), .ZN(new_n288));
  INV_X1    g087(.A(new_n283), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n290), .A2(G231gat), .A3(G233gat), .A4(new_n284), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n287), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n287), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n261), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n291), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n287), .A2(new_n291), .A3(new_n293), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n260), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G134gat), .B(G162gat), .Z(new_n303));
  NAND2_X1  g102(.A1(G85gat), .A2(G92gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT7), .B1(new_n304), .B2(KEYINPUT93), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(KEYINPUT93), .B2(new_n304), .ZN(new_n306));
  INV_X1    g105(.A(G99gat), .ZN(new_n307));
  INV_X1    g106(.A(G106gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT8), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(KEYINPUT93), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n311), .C1(G85gat), .C2(G92gat), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G99gat), .B(G106gat), .Z(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n227), .B2(new_n229), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT94), .ZN(new_n317));
  AND2_X1   g116(.A1(G232gat), .A2(G233gat), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n315), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n316), .A2(KEYINPUT94), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n303), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  INV_X1    g122(.A(new_n303), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n317), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n318), .A2(KEYINPUT41), .ZN(new_n327));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n325), .A3(new_n329), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n277), .B(new_n315), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n315), .A2(KEYINPUT10), .A3(new_n272), .A4(new_n276), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G230gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n334), .A2(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n341), .B1(new_n336), .B2(new_n337), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(new_n344), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n302), .A2(new_n333), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  AND2_X1   g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(G211gat), .A2(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G204gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n203), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n361), .A2(new_n362), .B1(KEYINPUT22), .B2(new_n357), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n364), .B2(KEYINPUT70), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  INV_X1    g165(.A(new_n359), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n257), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n371), .A2(KEYINPUT73), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  INV_X1    g176(.A(G141gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G148gat), .ZN(new_n379));
  INV_X1    g178(.A(G148gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G141gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n383));
  AND2_X1   g182(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n379), .A2(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G155gat), .B(G162gat), .Z(new_n386));
  AOI22_X1  g185(.A1(new_n376), .A2(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n375), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(G141gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(G148gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n386), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n356), .A2(new_n370), .B1(new_n388), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n387), .A2(new_n356), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n366), .B1(new_n365), .B2(new_n369), .ZN(new_n400));
  OAI211_X1 g199(.A(G228gat), .B(G233gat), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n366), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n365), .A2(new_n369), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n364), .B2(new_n367), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n364), .A2(new_n367), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n363), .A2(new_n408), .A3(new_n359), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n410), .B2(new_n366), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n404), .B(new_n405), .C1(new_n411), .C2(new_n387), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n401), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n401), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT31), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G50gat), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n414), .B2(new_n416), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424));
  INV_X1    g223(.A(G120gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G113gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(G113gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G127gat), .A2(G134gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(G127gat), .A2(G134gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT65), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n425), .B2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT65), .A3(G120gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n426), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G127gat), .ZN(new_n439));
  INV_X1    g238(.A(G134gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT1), .B1(new_n441), .B2(new_n430), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n429), .A2(new_n433), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT24), .ZN(new_n445));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(G169gat), .A2(G176gat), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n447), .A2(new_n448), .B1(KEYINPUT23), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G169gat), .ZN(new_n451));
  INV_X1    g250(.A(G176gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT23), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT64), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n455), .B2(new_n454), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n457), .A2(new_n458), .B1(new_n462), .B2(new_n450), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n449), .B(KEYINPUT26), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G183gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467));
  INV_X1    g266(.A(G190gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT28), .ZN(new_n471));
  AND4_X1   g270(.A1(new_n446), .A2(new_n465), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n443), .B1(new_n463), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n459), .A2(new_n464), .B1(new_n470), .B2(KEYINPUT28), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n469), .A2(new_n446), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n438), .A2(new_n442), .ZN(new_n477));
  XNOR2_X1  g276(.A(G113gat), .B(G120gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n433), .B1(new_n478), .B2(KEYINPUT1), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n450), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT25), .B1(new_n450), .B2(new_n456), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n476), .B(new_n480), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n473), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT33), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT67), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n487), .A2(KEYINPUT67), .A3(KEYINPUT32), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n490), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n487), .B2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n498), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n485), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n473), .A2(new_n484), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n485), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n485), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n496), .C1(new_n502), .C2(new_n503), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR4_X1   g316(.A1(new_n423), .A2(new_n514), .A3(new_n517), .A4(KEYINPUT35), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n520));
  XNOR2_X1  g319(.A(G1gat), .B(G29gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G57gat), .B(G85gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  AND3_X1   g323(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT74), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT74), .B1(new_n393), .B2(new_n394), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT3), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n443), .B1(new_n387), .B2(new_n356), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT75), .B1(new_n395), .B2(new_n480), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n387), .A2(new_n531), .A3(new_n443), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT4), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT4), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n395), .B2(new_n480), .ZN(new_n535));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT5), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n529), .A2(new_n533), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n480), .B1(new_n525), .B2(new_n526), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT76), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT76), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n480), .C1(new_n525), .C2(new_n526), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n530), .A2(new_n532), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n536), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n395), .A2(new_n480), .A3(KEYINPUT75), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n531), .B1(new_n387), .B2(new_n443), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n534), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n395), .A2(new_n480), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n537), .B1(new_n550), .B2(KEYINPUT4), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT5), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n524), .B(new_n539), .C1(new_n546), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n541), .A2(new_n543), .B1(new_n530), .B2(new_n532), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT5), .B(new_n552), .C1(new_n557), .C2(new_n536), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n524), .B1(new_n558), .B2(new_n539), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n519), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(KEYINPUT6), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n539), .B1(new_n546), .B2(new_n553), .ZN(new_n562));
  INV_X1    g361(.A(new_n524), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT81), .A3(new_n555), .A4(new_n554), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G64gat), .B(G92gat), .Z(new_n567));
  XNOR2_X1  g366(.A(G8gat), .B(G36gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G226gat), .A2(G233gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n457), .A2(new_n458), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n571), .A2(new_n481), .B1(new_n475), .B2(new_n474), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n572), .B2(KEYINPUT29), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n574));
  INV_X1    g373(.A(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n573), .A2(new_n403), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n403), .B1(new_n573), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n576), .ZN(new_n580));
  INV_X1    g379(.A(new_n403), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n403), .A3(new_n576), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n569), .B(KEYINPUT71), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n586), .A3(KEYINPUT30), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n569), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT82), .B1(new_n566), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n518), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n513), .A2(KEYINPUT68), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n504), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n496), .C1(new_n503), .C2(new_n502), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n597), .A2(new_n422), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n559), .B1(new_n556), .B2(KEYINPUT78), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n554), .A2(new_n601), .A3(new_n555), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n561), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n599), .B(new_n591), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n604), .B1(new_n600), .B2(new_n602), .ZN(new_n608));
  INV_X1    g407(.A(new_n591), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n423), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n514), .B2(new_n517), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT36), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n529), .A2(new_n533), .A3(new_n535), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n537), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n524), .B1(new_n616), .B2(KEYINPUT39), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n557), .A2(new_n536), .ZN(new_n618));
  INV_X1    g417(.A(new_n616), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n557), .A2(KEYINPUT80), .A3(new_n536), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n622), .A2(KEYINPUT39), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n617), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n609), .B1(new_n624), .B2(KEYINPUT40), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n623), .ZN(new_n627));
  INV_X1    g426(.A(new_n617), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n629), .B2(new_n564), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n422), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n569), .B1(new_n588), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT37), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n588), .A2(new_n633), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(new_n632), .A3(new_n635), .A4(new_n585), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n579), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n566), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n610), .B(new_n614), .C1(new_n631), .C2(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n255), .B(new_n355), .C1(new_n607), .C2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n608), .A2(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n608), .A2(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT96), .B(G1gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n609), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G8gat), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(G8gat), .B2(new_n649), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT98), .ZN(G1325gat));
  INV_X1    g458(.A(new_n614), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n642), .A2(G15gat), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n514), .A2(new_n517), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n642), .A2(new_n423), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n333), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n301), .A2(new_n671), .A3(new_n354), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  AOI21_X1  g472(.A(new_n255), .B1(new_n607), .B2(new_n641), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n645), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n675), .A2(G29gat), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT45), .Z(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n333), .B1(new_n607), .B2(new_n641), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT35), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n662), .A2(new_n686), .A3(new_n422), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n566), .A2(new_n591), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT82), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n591), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n608), .A2(new_n609), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n686), .B1(new_n693), .B2(new_n599), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n641), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n671), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n680), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n685), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n354), .A2(KEYINPUT101), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n354), .A2(KEYINPUT101), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n255), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n301), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n645), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G29gat), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT103), .B1(new_n706), .B2(new_n645), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n678), .B1(new_n708), .B2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n675), .A2(G36gat), .A3(new_n591), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n705), .B2(new_n591), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  AOI21_X1  g513(.A(new_n680), .B1(new_n696), .B2(new_n683), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n682), .A2(new_n681), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n660), .B(new_n704), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n662), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n675), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n718), .B2(KEYINPUT104), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n717), .A2(new_n725), .A3(G43gat), .ZN(new_n726));
  AOI211_X1 g525(.A(KEYINPUT105), .B(KEYINPUT47), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n614), .B(new_n703), .C1(new_n685), .C2(new_n697), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n726), .A3(new_n722), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n723), .B1(new_n727), .B2(new_n733), .ZN(G1330gat));
  NOR3_X1   g533(.A1(new_n675), .A2(G50gat), .A3(new_n422), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n706), .A2(new_n423), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(G50gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g537(.A1(new_n701), .A2(new_n702), .A3(new_n301), .A4(new_n671), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n695), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n645), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n268), .ZN(G1332gat));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n609), .B1(new_n743), .B2(new_n266), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n266), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n660), .ZN(new_n749));
  INV_X1    g548(.A(new_n662), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G71gat), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n749), .A2(G71gat), .B1(new_n740), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n423), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n301), .A2(new_n255), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n301), .B2(new_n255), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n353), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n685), .B2(new_n697), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n645), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G85gat), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT108), .B1(new_n762), .B2(new_n645), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n682), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n682), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n676), .A2(G85gat), .A3(new_n354), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n764), .A2(new_n765), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  OAI211_X1 g573(.A(new_n353), .B(new_n760), .C1(new_n715), .C2(new_n716), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n775), .B2(new_n591), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n701), .A2(G92gat), .A3(new_n591), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n768), .B2(new_n770), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(G92gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n762), .B2(new_n609), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT110), .B1(new_n784), .B2(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n786), .B(new_n789), .ZN(G1337gat));
  NAND2_X1  g589(.A1(new_n762), .A2(new_n660), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n792));
  OAI21_X1  g591(.A(G99gat), .B1(new_n791), .B2(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n662), .A2(new_n353), .A3(new_n307), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n792), .A2(new_n793), .B1(new_n772), .B2(new_n794), .ZN(G1338gat));
  OAI21_X1  g594(.A(G106gat), .B1(new_n775), .B2(new_n422), .ZN(new_n796));
  INV_X1    g595(.A(new_n701), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n308), .A3(new_n423), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT112), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n772), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n355), .A2(new_n702), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n240), .B1(new_n236), .B2(new_n238), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n244), .A2(new_n245), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n206), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n353), .A2(new_n253), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n353), .A2(new_n253), .A3(KEYINPUT114), .A4(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n336), .A2(new_n337), .A3(new_n341), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n343), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n349), .B1(new_n351), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n350), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n808), .B(new_n809), .C1(new_n818), .C2(new_n255), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n333), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n331), .A2(new_n253), .A3(new_n332), .A4(new_n805), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n822), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n817), .A2(new_n350), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n816), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n802), .B1(new_n828), .B2(new_n301), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n599), .A2(new_n591), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n645), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT115), .Z(new_n833));
  NAND2_X1  g632(.A1(new_n702), .A2(new_n436), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT116), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n829), .A2(new_n423), .A3(new_n750), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n591), .A3(new_n645), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n255), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1340gat));
  NAND3_X1  g639(.A1(new_n833), .A2(new_n425), .A3(new_n353), .ZN(new_n841));
  OAI21_X1  g640(.A(G120gat), .B1(new_n838), .B2(new_n701), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n439), .A3(new_n301), .ZN(new_n844));
  INV_X1    g643(.A(new_n832), .ZN(new_n845));
  AOI21_X1  g644(.A(G127gat), .B1(new_n845), .B2(new_n302), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n440), .A3(new_n671), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n838), .B2(new_n333), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n614), .A2(new_n423), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n591), .B1(new_n853), .B2(KEYINPUT118), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(KEYINPUT118), .B2(new_n853), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n302), .B1(new_n820), .B2(new_n827), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n645), .B(new_n855), .C1(new_n856), .C2(new_n802), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n378), .A3(new_n702), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n861), .B(new_n862), .C1(new_n255), .C2(new_n818), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n863), .A2(new_n333), .B1(new_n823), .B2(new_n826), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n864), .A2(new_n302), .B1(new_n702), .B2(new_n355), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n865), .B2(new_n423), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n860), .B(new_n423), .C1(new_n856), .C2(new_n802), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n676), .A2(new_n609), .A3(new_n660), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n866), .A2(new_n869), .A3(new_n255), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n859), .B1(new_n870), .B2(new_n378), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n380), .A3(new_n353), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT57), .B1(new_n829), .B2(new_n422), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n863), .A2(new_n333), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n824), .A2(new_n816), .A3(new_n825), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n302), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n860), .B(new_n423), .C1(new_n878), .C2(new_n802), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n353), .A3(new_n868), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n874), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n869), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n380), .C1(new_n883), .C2(new_n353), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n882), .B2(new_n884), .ZN(G1345gat));
  OR2_X1    g684(.A1(new_n866), .A2(new_n869), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n302), .A2(G155gat), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT119), .B1(new_n857), .B2(new_n301), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n257), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n301), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n886), .A2(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT120), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n886), .B2(new_n333), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n857), .A2(G162gat), .A3(new_n333), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n829), .A2(new_n645), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n599), .A2(new_n609), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n451), .A3(new_n702), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n645), .A2(new_n591), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n837), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n255), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n797), .A2(G176gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n452), .B1(new_n900), .B2(new_n354), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n904), .B2(new_n301), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n302), .A2(new_n466), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n900), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n916), .B(new_n920), .C1(new_n900), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n468), .A3(new_n671), .ZN(new_n923));
  OAI21_X1  g722(.A(G190gat), .B1(new_n904), .B2(new_n333), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n853), .A2(new_n591), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n897), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n203), .A3(new_n702), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n645), .A2(new_n591), .A3(new_n660), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n880), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(new_n702), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n934), .B2(new_n203), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n353), .A2(new_n360), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n929), .A2(KEYINPUT62), .A3(new_n936), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n880), .A2(new_n797), .A3(new_n932), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G204gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1353gat));
  OR3_X1    g741(.A1(new_n929), .A2(G211gat), .A3(new_n301), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n875), .A2(new_n879), .A3(new_n302), .A4(new_n932), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G211gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(KEYINPUT126), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT126), .B1(new_n945), .B2(new_n946), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(G218gat), .B1(new_n930), .B2(new_n671), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n671), .A2(G218gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n933), .B2(new_n954), .ZN(G1355gat));
endmodule


