

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717;

  XOR2_X1 U366 ( .A(n484), .B(n543), .Z(n599) );
  NOR2_X1 U367 ( .A1(n599), .A2(n600), .ZN(n517) );
  NAND2_X1 U368 ( .A1(n597), .A2(n596), .ZN(n600) );
  NOR2_X1 U369 ( .A1(n694), .A2(n582), .ZN(n406) );
  NOR2_X2 U370 ( .A1(n713), .A2(n399), .ZN(n533) );
  NOR2_X1 U371 ( .A1(n717), .A2(n716), .ZN(n373) );
  NOR2_X1 U372 ( .A1(n587), .A2(n557), .ZN(n555) );
  XNOR2_X1 U373 ( .A(n480), .B(n479), .ZN(n513) );
  NOR2_X1 U374 ( .A1(n560), .A2(n478), .ZN(n480) );
  AND2_X1 U375 ( .A1(n359), .A2(n348), .ZN(n623) );
  XNOR2_X1 U376 ( .A(n402), .B(KEYINPUT35), .ZN(n713) );
  NOR2_X1 U377 ( .A1(n522), .A2(n618), .ZN(n523) );
  NOR2_X1 U378 ( .A1(n513), .A2(n512), .ZN(n365) );
  XNOR2_X1 U379 ( .A(n360), .B(KEYINPUT19), .ZN(n560) );
  XNOR2_X1 U380 ( .A(n665), .B(n408), .ZN(n666) );
  XNOR2_X1 U381 ( .A(n498), .B(KEYINPUT4), .ZN(n462) );
  XNOR2_X1 U382 ( .A(KEYINPUT10), .B(n457), .ZN(n495) );
  XOR2_X1 U383 ( .A(G122), .B(G104), .Z(n488) );
  XOR2_X1 U384 ( .A(G110), .B(G119), .Z(n447) );
  XNOR2_X1 U385 ( .A(n365), .B(KEYINPUT22), .ZN(n531) );
  XNOR2_X1 U386 ( .A(n376), .B(KEYINPUT102), .ZN(n548) );
  OR2_X1 U387 ( .A1(n524), .A2(n525), .ZN(n376) );
  AND2_X1 U388 ( .A1(n662), .A2(n663), .ZN(n412) );
  XNOR2_X1 U389 ( .A(n547), .B(n375), .ZN(n587) );
  XNOR2_X1 U390 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n375) );
  NAND2_X1 U391 ( .A1(n393), .A2(n390), .ZN(n389) );
  NOR2_X1 U392 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U393 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U394 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n367) );
  XNOR2_X1 U395 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U396 ( .A1(n581), .A2(n412), .ZN(n707) );
  XNOR2_X1 U397 ( .A(n382), .B(n380), .ZN(n505) );
  XNOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n382) );
  NOR2_X1 U399 ( .A1(n381), .A2(G953), .ZN(n380) );
  INV_X1 U400 ( .A(G234), .ZN(n381) );
  XNOR2_X1 U401 ( .A(n495), .B(n427), .ZN(n701) );
  XNOR2_X1 U402 ( .A(G122), .B(KEYINPUT97), .ZN(n501) );
  XOR2_X1 U403 ( .A(G134), .B(KEYINPUT98), .Z(n502) );
  AND2_X1 U404 ( .A1(n581), .A2(n385), .ZN(n379) );
  INV_X1 U405 ( .A(n412), .ZN(n386) );
  XNOR2_X1 U406 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U407 ( .A1(n350), .A2(n354), .ZN(n574) );
  NOR2_X1 U408 ( .A1(n655), .A2(n407), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n384), .B(n383), .ZN(n511) );
  XNOR2_X1 U410 ( .A(KEYINPUT99), .B(G478), .ZN(n383) );
  OR2_X1 U411 ( .A1(n684), .A2(G902), .ZN(n384) );
  XNOR2_X1 U412 ( .A(n497), .B(n496), .ZN(n524) );
  NOR2_X1 U413 ( .A1(G902), .A2(n678), .ZN(n497) );
  NOR2_X1 U414 ( .A1(n689), .A2(G902), .ZN(n366) );
  XNOR2_X1 U415 ( .A(n510), .B(n353), .ZN(n568) );
  XNOR2_X1 U416 ( .A(KEYINPUT101), .B(KEYINPUT6), .ZN(n353) );
  OR2_X1 U417 ( .A1(G902), .A2(G237), .ZN(n472) );
  XOR2_X1 U418 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n422) );
  XOR2_X1 U419 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n442) );
  XNOR2_X1 U420 ( .A(n372), .B(n409), .ZN(n581) );
  NOR2_X1 U421 ( .A1(n567), .A2(n388), .ZN(n387) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n493) );
  XNOR2_X1 U423 ( .A(n462), .B(n413), .ZN(n702) );
  XNOR2_X1 U424 ( .A(G134), .B(G131), .ZN(n413) );
  XNOR2_X1 U425 ( .A(n461), .B(n358), .ZN(n463) );
  XNOR2_X1 U426 ( .A(n462), .B(n460), .ZN(n358) );
  NAND2_X1 U427 ( .A1(G237), .A2(G234), .ZN(n473) );
  INV_X1 U428 ( .A(KEYINPUT12), .ZN(n370) );
  XNOR2_X1 U429 ( .A(G131), .B(G140), .ZN(n490) );
  XNOR2_X1 U430 ( .A(n702), .B(G146), .ZN(n445) );
  XNOR2_X1 U431 ( .A(G107), .B(G104), .ZN(n414) );
  XOR2_X1 U432 ( .A(G110), .B(G101), .Z(n415) );
  XOR2_X1 U433 ( .A(G137), .B(G140), .Z(n426) );
  XNOR2_X1 U434 ( .A(n550), .B(n549), .ZN(n619) );
  NAND2_X1 U435 ( .A1(n590), .A2(n374), .ZN(n549) );
  NOR2_X1 U436 ( .A1(n587), .A2(n407), .ZN(n374) );
  NOR2_X1 U437 ( .A1(n389), .A2(n345), .ZN(n398) );
  XNOR2_X1 U438 ( .A(n397), .B(n351), .ZN(n396) );
  XNOR2_X1 U439 ( .A(n542), .B(n367), .ZN(n546) );
  XNOR2_X1 U440 ( .A(n434), .B(n433), .ZN(n689) );
  XNOR2_X1 U441 ( .A(n701), .B(n447), .ZN(n434) );
  XNOR2_X1 U442 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U443 ( .A(n346), .B(n508), .ZN(n684) );
  XNOR2_X1 U444 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U445 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n507) );
  XNOR2_X1 U446 ( .A(n371), .B(n368), .ZN(n678) );
  XNOR2_X1 U447 ( .A(n495), .B(n369), .ZN(n368) );
  XNOR2_X1 U448 ( .A(n492), .B(n489), .ZN(n371) );
  XNOR2_X1 U449 ( .A(n494), .B(n370), .ZN(n369) );
  NAND2_X1 U450 ( .A1(n585), .A2(n584), .ZN(n359) );
  XNOR2_X1 U451 ( .A(n404), .B(KEYINPUT75), .ZN(n585) );
  INV_X1 U452 ( .A(G953), .ZN(n709) );
  NOR2_X1 U453 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U454 ( .A1(n527), .A2(n529), .ZN(n528) );
  AND2_X1 U455 ( .A1(n600), .A2(KEYINPUT108), .ZN(n345) );
  XOR2_X1 U456 ( .A(n504), .B(n503), .Z(n346) );
  XOR2_X1 U457 ( .A(KEYINPUT5), .B(G119), .Z(n347) );
  XOR2_X1 U458 ( .A(n622), .B(KEYINPUT121), .Z(n348) );
  OR2_X1 U459 ( .A1(n707), .A2(n582), .ZN(n349) );
  AND2_X1 U460 ( .A1(n569), .A2(n568), .ZN(n350) );
  XNOR2_X1 U461 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n351) );
  INV_X1 U462 ( .A(n586), .ZN(n407) );
  XOR2_X1 U463 ( .A(n536), .B(KEYINPUT78), .Z(n352) );
  NAND2_X1 U464 ( .A1(n355), .A2(n387), .ZN(n372) );
  XNOR2_X1 U465 ( .A(n373), .B(KEYINPUT46), .ZN(n355) );
  XNOR2_X1 U466 ( .A(n364), .B(n471), .ZN(n579) );
  NOR2_X1 U467 ( .A1(n681), .A2(n691), .ZN(n361) );
  INV_X1 U468 ( .A(n356), .ZN(n547) );
  BUF_X1 U469 ( .A(n579), .Z(n356) );
  NOR2_X1 U470 ( .A1(n636), .A2(n691), .ZN(n638) );
  NAND2_X1 U471 ( .A1(n378), .A2(n628), .ZN(n362) );
  NAND2_X1 U472 ( .A1(n357), .A2(n455), .ZN(n459) );
  INV_X1 U473 ( .A(n456), .ZN(n357) );
  XNOR2_X1 U474 ( .A(n454), .B(n453), .ZN(n456) );
  NOR2_X1 U475 ( .A1(n579), .A2(n407), .ZN(n360) );
  NAND2_X1 U476 ( .A1(n694), .A2(n379), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n361), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U478 ( .A1(n668), .A2(n691), .ZN(n669) );
  XNOR2_X2 U479 ( .A(n362), .B(n629), .ZN(n631) );
  XNOR2_X2 U480 ( .A(n363), .B(n352), .ZN(n694) );
  NAND2_X1 U481 ( .A1(n535), .A2(n534), .ZN(n363) );
  XNOR2_X1 U482 ( .A(n521), .B(n520), .ZN(n618) );
  XNOR2_X2 U483 ( .A(n420), .B(G469), .ZN(n543) );
  NAND2_X1 U484 ( .A1(n664), .A2(n468), .ZN(n364) );
  NOR2_X1 U485 ( .A1(n685), .A2(n691), .ZN(n686) );
  XNOR2_X2 U486 ( .A(n366), .B(n435), .ZN(n597) );
  NOR2_X1 U487 ( .A1(n548), .A2(n587), .ZN(n593) );
  NAND2_X1 U488 ( .A1(n715), .A2(n377), .ZN(n399) );
  XNOR2_X1 U489 ( .A(n377), .B(G119), .ZN(G21) );
  XNOR2_X2 U490 ( .A(n400), .B(KEYINPUT32), .ZN(n377) );
  NOR2_X1 U491 ( .A1(n386), .A2(n468), .ZN(n385) );
  NOR2_X2 U492 ( .A1(G902), .A2(n632), .ZN(n446) );
  INV_X1 U493 ( .A(n661), .ZN(n388) );
  NOR2_X1 U494 ( .A1(n600), .A2(n543), .ZN(n553) );
  INV_X1 U495 ( .A(n554), .ZN(n391) );
  AND2_X1 U496 ( .A1(n543), .A2(KEYINPUT108), .ZN(n392) );
  NOR2_X1 U497 ( .A1(n543), .A2(KEYINPUT108), .ZN(n394) );
  INV_X1 U498 ( .A(n600), .ZN(n395) );
  NAND2_X1 U499 ( .A1(n398), .A2(n396), .ZN(n557) );
  NAND2_X1 U500 ( .A1(n552), .A2(n586), .ZN(n397) );
  NAND2_X1 U501 ( .A1(n531), .A2(n528), .ZN(n400) );
  XNOR2_X2 U502 ( .A(n401), .B(KEYINPUT104), .ZN(n715) );
  NAND2_X1 U503 ( .A1(n531), .A2(n532), .ZN(n401) );
  NAND2_X1 U504 ( .A1(n403), .A2(n526), .ZN(n402) );
  XNOR2_X1 U505 ( .A(n523), .B(KEYINPUT34), .ZN(n403) );
  NAND2_X1 U506 ( .A1(n405), .A2(n349), .ZN(n404) );
  XNOR2_X1 U507 ( .A(n406), .B(KEYINPUT77), .ZN(n405) );
  BUF_X1 U508 ( .A(n682), .Z(n687) );
  XNOR2_X1 U509 ( .A(n605), .B(KEYINPUT103), .ZN(n552) );
  INV_X1 U510 ( .A(n605), .ZN(n510) );
  XNOR2_X2 U511 ( .A(n438), .B(KEYINPUT3), .ZN(n448) );
  XNOR2_X2 U512 ( .A(G101), .B(G113), .ZN(n438) );
  XNOR2_X1 U513 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n408) );
  XNOR2_X1 U514 ( .A(KEYINPUT48), .B(KEYINPUT69), .ZN(n409) );
  XOR2_X1 U515 ( .A(n444), .B(n443), .Z(n410) );
  XOR2_X1 U516 ( .A(KEYINPUT53), .B(n624), .Z(G75) );
  INV_X1 U517 ( .A(KEYINPUT33), .ZN(n518) );
  XNOR2_X1 U518 ( .A(n445), .B(n410), .ZN(n632) );
  INV_X1 U519 ( .A(n426), .ZN(n427) );
  INV_X1 U520 ( .A(n630), .ZN(n584) );
  XNOR2_X1 U521 ( .A(n632), .B(n633), .ZN(n634) );
  XNOR2_X1 U522 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U523 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U524 ( .A(KEYINPUT82), .B(n625), .ZN(n691) );
  XNOR2_X2 U525 ( .A(G143), .B(G128), .ZN(n498) );
  XNOR2_X1 U526 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U527 ( .A(n426), .B(n416), .Z(n418) );
  NAND2_X1 U528 ( .A1(G227), .A2(n709), .ZN(n417) );
  XNOR2_X1 U529 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U530 ( .A(n445), .B(n419), .ZN(n673) );
  NOR2_X1 U531 ( .A1(n673), .A2(G902), .ZN(n420) );
  XOR2_X1 U532 ( .A(KEYINPUT73), .B(KEYINPUT25), .Z(n424) );
  XOR2_X1 U533 ( .A(G902), .B(KEYINPUT15), .Z(n626) );
  INV_X1 U534 ( .A(n626), .ZN(n468) );
  NAND2_X1 U535 ( .A1(G234), .A2(n468), .ZN(n421) );
  XNOR2_X1 U536 ( .A(n422), .B(n421), .ZN(n436) );
  NAND2_X1 U537 ( .A1(n436), .A2(G217), .ZN(n423) );
  XNOR2_X1 U538 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U539 ( .A(KEYINPUT90), .B(n425), .ZN(n435) );
  XNOR2_X2 U540 ( .A(G146), .B(G125), .ZN(n457) );
  XOR2_X1 U541 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U542 ( .A(G128), .B(KEYINPUT88), .ZN(n428) );
  XNOR2_X1 U543 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U544 ( .A(n430), .B(KEYINPUT24), .Z(n432) );
  NAND2_X1 U545 ( .A1(G221), .A2(n505), .ZN(n431) );
  NAND2_X1 U546 ( .A1(G221), .A2(n436), .ZN(n437) );
  XOR2_X1 U547 ( .A(KEYINPUT21), .B(n437), .Z(n596) );
  XNOR2_X1 U548 ( .A(G116), .B(G137), .ZN(n439) );
  XNOR2_X1 U549 ( .A(n347), .B(n439), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n448), .B(n440), .ZN(n444) );
  NAND2_X1 U551 ( .A1(n493), .A2(G210), .ZN(n441) );
  XNOR2_X1 U552 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X2 U553 ( .A(n446), .B(G472), .ZN(n605) );
  XOR2_X1 U554 ( .A(n488), .B(n447), .Z(n450) );
  XOR2_X1 U555 ( .A(G116), .B(G107), .Z(n500) );
  XNOR2_X1 U556 ( .A(n448), .B(n500), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n449), .B(n450), .ZN(n452) );
  XOR2_X1 U558 ( .A(KEYINPUT70), .B(KEYINPUT16), .Z(n451) );
  XNOR2_X1 U559 ( .A(n452), .B(n451), .ZN(n697) );
  INV_X1 U560 ( .A(n457), .ZN(n455) );
  XOR2_X1 U561 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n454) );
  XNOR2_X1 U562 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n453) );
  NAND2_X1 U563 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U564 ( .A1(n459), .A2(n458), .ZN(n461) );
  NAND2_X1 U565 ( .A1(G224), .A2(n709), .ZN(n460) );
  NAND2_X1 U566 ( .A1(n697), .A2(n463), .ZN(n467) );
  INV_X1 U567 ( .A(n463), .ZN(n465) );
  INV_X1 U568 ( .A(n697), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U570 ( .A1(n467), .A2(n466), .ZN(n664) );
  NAND2_X1 U571 ( .A1(G210), .A2(n472), .ZN(n470) );
  INV_X1 U572 ( .A(KEYINPUT85), .ZN(n469) );
  NAND2_X1 U573 ( .A1(G214), .A2(n472), .ZN(n586) );
  XNOR2_X1 U574 ( .A(n473), .B(KEYINPUT14), .ZN(n474) );
  NAND2_X1 U575 ( .A1(G952), .A2(n474), .ZN(n617) );
  NOR2_X1 U576 ( .A1(G953), .A2(n617), .ZN(n539) );
  NAND2_X1 U577 ( .A1(G902), .A2(n474), .ZN(n475) );
  XOR2_X1 U578 ( .A(KEYINPUT86), .B(n475), .Z(n476) );
  NAND2_X1 U579 ( .A1(G953), .A2(n476), .ZN(n537) );
  NOR2_X1 U580 ( .A1(G898), .A2(n537), .ZN(n477) );
  NOR2_X1 U581 ( .A1(n539), .A2(n477), .ZN(n478) );
  XNOR2_X1 U582 ( .A(KEYINPUT79), .B(KEYINPUT0), .ZN(n479) );
  INV_X1 U583 ( .A(KEYINPUT87), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n513), .B(n481), .ZN(n522) );
  NOR2_X1 U585 ( .A1(n510), .A2(n522), .ZN(n482) );
  NAND2_X1 U586 ( .A1(n553), .A2(n482), .ZN(n483) );
  XNOR2_X1 U587 ( .A(KEYINPUT94), .B(n483), .ZN(n642) );
  XNOR2_X1 U588 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n484) );
  NAND2_X1 U589 ( .A1(n510), .A2(n517), .ZN(n607) );
  NOR2_X1 U590 ( .A1(n513), .A2(n607), .ZN(n486) );
  XNOR2_X1 U591 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U593 ( .A(KEYINPUT95), .B(n487), .Z(n658) );
  NAND2_X1 U594 ( .A1(n642), .A2(n658), .ZN(n509) );
  XNOR2_X1 U595 ( .A(G143), .B(n488), .ZN(n489) );
  XOR2_X1 U596 ( .A(KEYINPUT11), .B(G113), .Z(n491) );
  XNOR2_X1 U597 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U598 ( .A1(n493), .A2(G214), .ZN(n494) );
  XNOR2_X1 U599 ( .A(KEYINPUT13), .B(G475), .ZN(n496) );
  INV_X1 U600 ( .A(n498), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n500), .B(n499), .ZN(n504) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U603 ( .A1(G217), .A2(n505), .ZN(n506) );
  NOR2_X1 U604 ( .A1(n524), .A2(n511), .ZN(n647) );
  XNOR2_X1 U605 ( .A(KEYINPUT100), .B(n647), .ZN(n572) );
  NAND2_X1 U606 ( .A1(n524), .A2(n511), .ZN(n655) );
  INV_X1 U607 ( .A(n655), .ZN(n652) );
  NOR2_X1 U608 ( .A1(n572), .A2(n652), .ZN(n588) );
  INV_X1 U609 ( .A(n588), .ZN(n562) );
  NAND2_X1 U610 ( .A1(n509), .A2(n562), .ZN(n516) );
  INV_X1 U611 ( .A(n511), .ZN(n525) );
  INV_X1 U612 ( .A(n548), .ZN(n590) );
  NAND2_X1 U613 ( .A1(n590), .A2(n596), .ZN(n512) );
  NAND2_X1 U614 ( .A1(n597), .A2(n531), .ZN(n514) );
  NOR2_X1 U615 ( .A1(n568), .A2(n514), .ZN(n515) );
  NAND2_X1 U616 ( .A1(n599), .A2(n515), .ZN(n639) );
  AND2_X1 U617 ( .A1(n516), .A2(n639), .ZN(n535) );
  NAND2_X1 U618 ( .A1(n517), .A2(n568), .ZN(n521) );
  XOR2_X1 U619 ( .A(KEYINPUT80), .B(KEYINPUT105), .Z(n519) );
  NAND2_X1 U620 ( .A1(n525), .A2(n524), .ZN(n559) );
  INV_X1 U621 ( .A(n559), .ZN(n526) );
  NOR2_X1 U622 ( .A1(n599), .A2(n568), .ZN(n527) );
  INV_X1 U623 ( .A(n597), .ZN(n529) );
  INV_X1 U624 ( .A(n599), .ZN(n576) );
  NOR2_X1 U625 ( .A1(n576), .A2(n552), .ZN(n530) );
  AND2_X1 U626 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  INV_X1 U628 ( .A(KEYINPUT45), .ZN(n536) );
  XNOR2_X1 U629 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n582) );
  NOR2_X1 U630 ( .A1(G900), .A2(n537), .ZN(n538) );
  NOR2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U632 ( .A(KEYINPUT74), .B(n540), .Z(n554) );
  NAND2_X1 U633 ( .A1(n554), .A2(n596), .ZN(n541) );
  NOR2_X1 U634 ( .A1(n597), .A2(n541), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n552), .A2(n569), .ZN(n542) );
  INV_X1 U636 ( .A(n543), .ZN(n544) );
  XNOR2_X1 U637 ( .A(n544), .B(KEYINPUT110), .ZN(n545) );
  NAND2_X1 U638 ( .A1(n546), .A2(n545), .ZN(n561) );
  XOR2_X1 U639 ( .A(KEYINPUT112), .B(KEYINPUT41), .Z(n550) );
  NOR2_X1 U640 ( .A1(n561), .A2(n619), .ZN(n551) );
  XNOR2_X1 U641 ( .A(n551), .B(KEYINPUT42), .ZN(n717) );
  XOR2_X1 U642 ( .A(n555), .B(KEYINPUT39), .Z(n573) );
  AND2_X1 U643 ( .A1(n652), .A2(n573), .ZN(n556) );
  XNOR2_X1 U644 ( .A(KEYINPUT40), .B(n556), .ZN(n716) );
  OR2_X1 U645 ( .A1(n356), .A2(n557), .ZN(n558) );
  NOR2_X1 U646 ( .A1(n559), .A2(n558), .ZN(n650) );
  NOR2_X2 U647 ( .A1(n561), .A2(n560), .ZN(n651) );
  NAND2_X1 U648 ( .A1(n651), .A2(n562), .ZN(n563) );
  NOR2_X1 U649 ( .A1(KEYINPUT67), .A2(n563), .ZN(n564) );
  XOR2_X1 U650 ( .A(KEYINPUT47), .B(n564), .Z(n565) );
  NOR2_X1 U651 ( .A1(n650), .A2(n565), .ZN(n566) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(n566), .ZN(n567) );
  NOR2_X1 U653 ( .A1(n356), .A2(n574), .ZN(n570) );
  XNOR2_X1 U654 ( .A(KEYINPUT36), .B(n570), .ZN(n571) );
  NAND2_X1 U655 ( .A1(n571), .A2(n576), .ZN(n661) );
  NAND2_X1 U656 ( .A1(n573), .A2(n572), .ZN(n662) );
  XNOR2_X1 U657 ( .A(n574), .B(KEYINPUT106), .ZN(n575) );
  XNOR2_X1 U658 ( .A(KEYINPUT43), .B(n577), .ZN(n578) );
  XNOR2_X1 U659 ( .A(n578), .B(KEYINPUT107), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n580), .A2(n356), .ZN(n663) );
  AND2_X1 U661 ( .A1(n694), .A2(n707), .ZN(n583) );
  AND2_X1 U662 ( .A1(KEYINPUT2), .A2(n583), .ZN(n630) );
  NOR2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U665 ( .A1(n407), .A2(n591), .ZN(n592) );
  NOR2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n618), .A2(n594), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT120), .ZN(n614) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT49), .B(n598), .Z(n604) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT117), .ZN(n602) );
  XNOR2_X1 U673 ( .A(KEYINPUT50), .B(n602), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n611) );
  XOR2_X1 U677 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n609) );
  XNOR2_X1 U678 ( .A(KEYINPUT51), .B(n609), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n612), .A2(n619), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U682 ( .A(n615), .B(KEYINPUT52), .ZN(n616) );
  NOR2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n621) );
  NOR2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U685 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U686 ( .A1(n709), .A2(n623), .ZN(n624) );
  NOR2_X1 U687 ( .A1(G952), .A2(n709), .ZN(n625) );
  INV_X1 U688 ( .A(KEYINPUT64), .ZN(n629) );
  NAND2_X1 U689 ( .A1(KEYINPUT2), .A2(n626), .ZN(n627) );
  XNOR2_X1 U690 ( .A(n627), .B(KEYINPUT66), .ZN(n628) );
  NOR2_X4 U691 ( .A1(n631), .A2(n630), .ZN(n682) );
  NAND2_X1 U692 ( .A1(n682), .A2(G472), .ZN(n635) );
  XOR2_X1 U693 ( .A(KEYINPUT62), .B(KEYINPUT81), .Z(n633) );
  XNOR2_X1 U694 ( .A(KEYINPUT63), .B(KEYINPUT113), .ZN(n637) );
  XNOR2_X1 U695 ( .A(n638), .B(n637), .ZN(G57) );
  XNOR2_X1 U696 ( .A(G101), .B(n639), .ZN(G3) );
  NOR2_X1 U697 ( .A1(n642), .A2(n655), .ZN(n640) );
  XOR2_X1 U698 ( .A(KEYINPUT114), .B(n640), .Z(n641) );
  XNOR2_X1 U699 ( .A(G104), .B(n641), .ZN(G6) );
  INV_X1 U700 ( .A(n647), .ZN(n657) );
  NOR2_X1 U701 ( .A1(n657), .A2(n642), .ZN(n646) );
  XOR2_X1 U702 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n644) );
  XNOR2_X1 U703 ( .A(G107), .B(KEYINPUT27), .ZN(n643) );
  XNOR2_X1 U704 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U705 ( .A(n646), .B(n645), .ZN(G9) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U707 ( .A1(n647), .A2(n651), .ZN(n648) );
  XNOR2_X1 U708 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U709 ( .A(G143), .B(n650), .Z(G45) );
  XNOR2_X1 U710 ( .A(G146), .B(KEYINPUT116), .ZN(n654) );
  NAND2_X1 U711 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U712 ( .A(n654), .B(n653), .ZN(G48) );
  NOR2_X1 U713 ( .A1(n658), .A2(n655), .ZN(n656) );
  XOR2_X1 U714 ( .A(G113), .B(n656), .Z(G15) );
  NOR2_X1 U715 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U716 ( .A(G116), .B(n659), .Z(G18) );
  XOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .Z(n660) );
  XNOR2_X1 U718 ( .A(n661), .B(n660), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n662), .ZN(G36) );
  XNOR2_X1 U720 ( .A(G140), .B(n663), .ZN(G42) );
  NAND2_X1 U721 ( .A1(n682), .A2(G210), .ZN(n667) );
  BUF_X1 U722 ( .A(n664), .Z(n665) );
  XNOR2_X1 U723 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U724 ( .A(KEYINPUT56), .B(n669), .ZN(G51) );
  XOR2_X1 U725 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n671) );
  XNOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U728 ( .A(n673), .B(n672), .Z(n675) );
  NAND2_X1 U729 ( .A1(n687), .A2(G469), .ZN(n674) );
  XNOR2_X1 U730 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U731 ( .A1(n676), .A2(n691), .ZN(G54) );
  NAND2_X1 U732 ( .A1(n682), .A2(G475), .ZN(n680) );
  INV_X1 U733 ( .A(KEYINPUT59), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U735 ( .A1(G478), .A2(n682), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n683), .B(n684), .ZN(n685) );
  XNOR2_X1 U737 ( .A(KEYINPUT124), .B(n686), .ZN(G63) );
  NAND2_X1 U738 ( .A1(G217), .A2(n687), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U740 ( .A1(n691), .A2(n690), .ZN(G66) );
  NAND2_X1 U741 ( .A1(G953), .A2(G224), .ZN(n692) );
  XNOR2_X1 U742 ( .A(KEYINPUT61), .B(n692), .ZN(n693) );
  NAND2_X1 U743 ( .A1(n693), .A2(G898), .ZN(n696) );
  NAND2_X1 U744 ( .A1(n694), .A2(n709), .ZN(n695) );
  NAND2_X1 U745 ( .A1(n696), .A2(n695), .ZN(n700) );
  OR2_X1 U746 ( .A1(n709), .A2(G898), .ZN(n698) );
  NAND2_X1 U747 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U748 ( .A(n700), .B(n699), .Z(G69) );
  XNOR2_X1 U749 ( .A(n702), .B(n701), .ZN(n703) );
  XOR2_X1 U750 ( .A(n703), .B(KEYINPUT125), .Z(n708) );
  XOR2_X1 U751 ( .A(G227), .B(n708), .Z(n704) );
  NAND2_X1 U752 ( .A1(n704), .A2(G900), .ZN(n705) );
  NAND2_X1 U753 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U754 ( .A(n706), .B(KEYINPUT126), .ZN(n712) );
  XNOR2_X1 U755 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U756 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U757 ( .A1(n712), .A2(n711), .ZN(G72) );
  XNOR2_X1 U758 ( .A(n713), .B(G122), .ZN(n714) );
  XNOR2_X1 U759 ( .A(n714), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U760 ( .A(G110), .B(n715), .ZN(G12) );
  XOR2_X1 U761 ( .A(G131), .B(n716), .Z(G33) );
  XOR2_X1 U762 ( .A(G137), .B(n717), .Z(G39) );
endmodule

