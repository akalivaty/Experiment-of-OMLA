

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n658), .A2(n551), .ZN(n642) );
  NOR2_X2 U557 ( .A1(n724), .A2(n738), .ZN(n725) );
  BUF_X1 U558 ( .A(n568), .Z(n523) );
  NOR2_X1 U559 ( .A1(G2104), .A2(n531), .ZN(n568) );
  XNOR2_X1 U560 ( .A(KEYINPUT64), .B(n694), .ZN(n701) );
  AND2_X1 U561 ( .A1(n690), .A2(n689), .ZN(n691) );
  BUF_X1 U562 ( .A(n571), .Z(n537) );
  XNOR2_X1 U563 ( .A(n732), .B(KEYINPUT99), .ZN(n733) );
  XNOR2_X1 U564 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n751) );
  INV_X1 U565 ( .A(n985), .ZN(n757) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  INV_X1 U567 ( .A(n695), .ZN(n742) );
  AND2_X1 U568 ( .A1(n827), .A2(n817), .ZN(n524) );
  NAND2_X1 U569 ( .A1(n762), .A2(n756), .ZN(n525) );
  NOR2_X1 U570 ( .A1(n714), .A2(n713), .ZN(n700) );
  INV_X1 U571 ( .A(KEYINPUT31), .ZN(n732) );
  XNOR2_X1 U572 ( .A(n734), .B(n733), .ZN(n735) );
  INV_X1 U573 ( .A(KEYINPUT101), .ZN(n748) );
  XNOR2_X1 U574 ( .A(n752), .B(n751), .ZN(n753) );
  NAND2_X1 U575 ( .A1(n764), .A2(n774), .ZN(n765) );
  INV_X1 U576 ( .A(KEYINPUT74), .ZN(n581) );
  XNOR2_X1 U577 ( .A(n581), .B(KEYINPUT13), .ZN(n582) );
  XNOR2_X1 U578 ( .A(n583), .B(n582), .ZN(n584) );
  INV_X1 U579 ( .A(KEYINPUT17), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n524), .A2(n818), .ZN(n819) );
  NOR2_X1 U581 ( .A1(n658), .A2(G651), .ZN(n652) );
  NAND2_X1 U582 ( .A1(n889), .A2(G137), .ZN(n690) );
  NAND2_X1 U583 ( .A1(n588), .A2(n587), .ZN(n987) );
  NAND2_X1 U584 ( .A1(n531), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U585 ( .A(n526), .B(KEYINPUT65), .ZN(n571) );
  NAND2_X1 U586 ( .A1(G102), .A2(n571), .ZN(n530) );
  XNOR2_X2 U587 ( .A(n528), .B(n527), .ZN(n889) );
  NAND2_X1 U588 ( .A1(G138), .A2(n889), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n535) );
  INV_X1 U590 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U591 ( .A1(G126), .A2(n523), .ZN(n533) );
  AND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U593 ( .A1(G114), .A2(n895), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U595 ( .A1(n535), .A2(n534), .ZN(G164) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U597 ( .A1(G123), .A2(n523), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(KEYINPUT18), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G99), .A2(n537), .ZN(n539) );
  NAND2_X1 U600 ( .A1(G111), .A2(n895), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G135), .A2(n889), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT79), .B(n540), .ZN(n541) );
  NOR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n929) );
  XNOR2_X1 U606 ( .A(G2096), .B(n929), .ZN(n545) );
  OR2_X1 U607 ( .A1(G2100), .A2(n545), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NOR2_X1 U611 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U612 ( .A1(n644), .A2(G89), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT4), .B(n546), .ZN(n549) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n658) );
  INV_X1 U615 ( .A(G651), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n642), .A2(G76), .ZN(n547) );
  XOR2_X1 U617 ( .A(KEYINPUT77), .B(n547), .Z(n548) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(n550), .ZN(n559) );
  NOR2_X1 U620 ( .A1(G543), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n657) );
  NAND2_X1 U623 ( .A1(G63), .A2(n657), .ZN(n555) );
  NAND2_X1 U624 ( .A1(G51), .A2(n652), .ZN(n554) );
  NAND2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n557) );
  XOR2_X1 U626 ( .A(KEYINPUT78), .B(KEYINPUT6), .Z(n556) );
  XNOR2_X1 U627 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  NAND2_X1 U630 ( .A1(G88), .A2(n644), .ZN(n562) );
  NAND2_X1 U631 ( .A1(G75), .A2(n642), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U633 ( .A(KEYINPUT84), .B(n563), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G62), .A2(n657), .ZN(n565) );
  NAND2_X1 U635 ( .A1(G50), .A2(n652), .ZN(n564) );
  NAND2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U637 ( .A1(n567), .A2(n566), .ZN(G166) );
  INV_X1 U638 ( .A(G166), .ZN(G303) );
  NAND2_X1 U639 ( .A1(G125), .A2(n568), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G113), .A2(n895), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n687) );
  NAND2_X1 U642 ( .A1(G101), .A2(n571), .ZN(n572) );
  XOR2_X1 U643 ( .A(KEYINPUT23), .B(n572), .Z(n692) );
  NAND2_X1 U644 ( .A1(n692), .A2(n690), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n687), .A2(n573), .ZN(G160) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n837) );
  NAND2_X1 U649 ( .A1(n837), .A2(G567), .ZN(n575) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U651 ( .A1(n657), .A2(G56), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n576), .B(KEYINPUT14), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n642), .A2(G68), .ZN(n577) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(n577), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n644), .A2(G81), .ZN(n578) );
  XOR2_X1 U656 ( .A(n578), .B(KEYINPUT12), .Z(n579) );
  NOR2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT75), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G43), .A2(n652), .ZN(n587) );
  INV_X1 U661 ( .A(G860), .ZN(n618) );
  OR2_X1 U662 ( .A1(n987), .A2(n618), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G52), .A2(n652), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n657), .A2(G64), .ZN(n589) );
  XNOR2_X1 U665 ( .A(KEYINPUT69), .B(n589), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G90), .A2(n644), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G77), .A2(n642), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U669 ( .A(KEYINPUT70), .B(n592), .Z(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT9), .B(n593), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT71), .ZN(G171) );
  INV_X1 U674 ( .A(G171), .ZN(G301) );
  NAND2_X1 U675 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G66), .A2(n657), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G79), .A2(n642), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G92), .A2(n644), .ZN(n602) );
  NAND2_X1 U680 ( .A1(G54), .A2(n652), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n606), .B(n605), .ZN(n906) );
  INV_X1 U685 ( .A(G868), .ZN(n671) );
  NAND2_X1 U686 ( .A1(n906), .A2(n671), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U688 ( .A1(G91), .A2(n644), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G65), .A2(n657), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n642), .A2(G78), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT72), .B(n611), .Z(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n652), .A2(G53), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G299) );
  XOR2_X1 U696 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U698 ( .A1(G286), .A2(n671), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(G297) );
  NAND2_X1 U700 ( .A1(n618), .A2(G559), .ZN(n619) );
  INV_X1 U701 ( .A(n906), .ZN(n990) );
  NAND2_X1 U702 ( .A1(n619), .A2(n990), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(G868), .A2(n987), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n990), .A2(G868), .ZN(n621) );
  NOR2_X1 U706 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G67), .A2(n657), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G80), .A2(n642), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G93), .A2(n644), .ZN(n627) );
  NAND2_X1 U712 ( .A1(G55), .A2(n652), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n670) );
  XNOR2_X1 U715 ( .A(n987), .B(KEYINPUT80), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n990), .A2(G559), .ZN(n630) );
  XNOR2_X1 U717 ( .A(n631), .B(n630), .ZN(n667) );
  XOR2_X1 U718 ( .A(n667), .B(KEYINPUT81), .Z(n632) );
  NOR2_X1 U719 ( .A1(G860), .A2(n632), .ZN(n633) );
  XOR2_X1 U720 ( .A(n670), .B(n633), .Z(G145) );
  NAND2_X1 U721 ( .A1(n642), .A2(G72), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n652), .A2(G47), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n657), .A2(G60), .ZN(n634) );
  NAND2_X1 U724 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U725 ( .A1(G85), .A2(n644), .ZN(n636) );
  XOR2_X1 U726 ( .A(KEYINPUT66), .B(n636), .Z(n637) );
  NOR2_X1 U727 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n641), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U730 ( .A1(G73), .A2(n642), .ZN(n643) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n643), .Z(n649) );
  NAND2_X1 U732 ( .A1(G86), .A2(n644), .ZN(n646) );
  NAND2_X1 U733 ( .A1(G61), .A2(n657), .ZN(n645) );
  NAND2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U735 ( .A(KEYINPUT83), .B(n647), .Z(n648) );
  NOR2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(G48), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G49), .A2(n652), .ZN(n654) );
  NAND2_X1 U740 ( .A1(G74), .A2(G651), .ZN(n653) );
  NAND2_X1 U741 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U742 ( .A(KEYINPUT82), .B(n655), .ZN(n656) );
  NOR2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n658), .A2(G87), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(G288) );
  XOR2_X1 U746 ( .A(n670), .B(KEYINPUT85), .Z(n661) );
  XNOR2_X1 U747 ( .A(n661), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U748 ( .A(G290), .B(G305), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n662), .B(G303), .ZN(n663) );
  XNOR2_X1 U750 ( .A(n664), .B(n663), .ZN(n666) );
  INV_X1 U751 ( .A(G299), .ZN(n713) );
  XNOR2_X1 U752 ( .A(G288), .B(n713), .ZN(n665) );
  XNOR2_X1 U753 ( .A(n666), .B(n665), .ZN(n905) );
  XNOR2_X1 U754 ( .A(n905), .B(n667), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n668), .A2(G868), .ZN(n669) );
  XNOR2_X1 U756 ( .A(n669), .B(KEYINPUT86), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n675), .ZN(n677) );
  XOR2_X1 U762 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n676) );
  XNOR2_X1 U763 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U764 ( .A1(G2072), .A2(n678), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U768 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G96), .A2(n681), .ZN(n926) );
  NAND2_X1 U770 ( .A1(n926), .A2(G2106), .ZN(n685) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U772 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U773 ( .A1(G108), .A2(n683), .ZN(n925) );
  NAND2_X1 U774 ( .A1(n925), .A2(G567), .ZN(n684) );
  NAND2_X1 U775 ( .A1(n685), .A2(n684), .ZN(n842) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n842), .A2(n686), .ZN(n841) );
  NAND2_X1 U778 ( .A1(n841), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G40), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n794) );
  XNOR2_X1 U782 ( .A(n794), .B(KEYINPUT95), .ZN(n693) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n795) );
  NAND2_X1 U784 ( .A1(n693), .A2(n795), .ZN(n694) );
  INV_X1 U785 ( .A(n701), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n742), .A2(G2084), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n724), .A2(G8), .ZN(n740) );
  NAND2_X1 U788 ( .A1(G8), .A2(n701), .ZN(n779) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n779), .ZN(n738) );
  NAND2_X1 U790 ( .A1(G2072), .A2(n695), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U792 ( .A(G1956), .ZN(n1014) );
  NOR2_X1 U793 ( .A1(n695), .A2(n1014), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n714) );
  XNOR2_X1 U795 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n699) );
  XNOR2_X1 U796 ( .A(n700), .B(n699), .ZN(n718) );
  INV_X1 U797 ( .A(G1996), .ZN(n959) );
  NOR2_X1 U798 ( .A1(n701), .A2(n959), .ZN(n702) );
  XOR2_X1 U799 ( .A(n702), .B(KEYINPUT26), .Z(n704) );
  NAND2_X1 U800 ( .A1(n742), .A2(G1341), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U802 ( .A1(n987), .A2(n705), .ZN(n706) );
  OR2_X1 U803 ( .A1(n706), .A2(n990), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n990), .A2(n706), .ZN(n710) );
  NAND2_X1 U805 ( .A1(G2067), .A2(n695), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n742), .A2(G1348), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n719), .B(KEYINPUT29), .ZN(n723) );
  XOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .Z(n965) );
  NAND2_X1 U815 ( .A1(n965), .A2(n695), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n742), .A2(G1961), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n729) );
  NOR2_X1 U818 ( .A1(G301), .A2(n729), .ZN(n722) );
  NOR2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n736) );
  XNOR2_X1 U820 ( .A(KEYINPUT98), .B(n725), .ZN(n726) );
  NAND2_X1 U821 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U822 ( .A(n727), .B(KEYINPUT30), .ZN(n728) );
  NOR2_X1 U823 ( .A1(G168), .A2(n728), .ZN(n731) );
  AND2_X1 U824 ( .A1(G301), .A2(n729), .ZN(n730) );
  NOR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n734) );
  OR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U827 ( .A(KEYINPUT100), .B(n741), .Z(n737) );
  NOR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n754) );
  NAND2_X1 U830 ( .A1(n741), .A2(G286), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n742), .A2(G2090), .ZN(n744) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n779), .ZN(n743) );
  NOR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n745), .A2(G303), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(G8), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n762) );
  NOR2_X1 U839 ( .A1(G303), .A2(G1971), .ZN(n755) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NOR2_X1 U841 ( .A1(n755), .A2(n980), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NOR2_X1 U843 ( .A1(n779), .A2(n757), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n525), .A2(n758), .ZN(n759) );
  NOR2_X1 U845 ( .A1(KEYINPUT103), .A2(n759), .ZN(n766) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n763), .A2(n779), .ZN(n774) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n776) );
  INV_X1 U852 ( .A(KEYINPUT103), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n980), .A2(KEYINPUT33), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n980), .A2(KEYINPUT103), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U857 ( .A1(n779), .A2(n771), .ZN(n772) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n998) );
  NAND2_X1 U859 ( .A1(n772), .A2(n998), .ZN(n773) );
  AND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n782) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U863 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(n780), .B(KEYINPUT96), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n820) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n829) );
  NAND2_X1 U868 ( .A1(G128), .A2(n523), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G116), .A2(n895), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n785), .Z(n792) );
  NAND2_X1 U872 ( .A1(n889), .A2(G140), .ZN(n786) );
  XNOR2_X1 U873 ( .A(KEYINPUT89), .B(n786), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n537), .A2(G104), .ZN(n787) );
  XOR2_X1 U875 ( .A(KEYINPUT88), .B(n787), .Z(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U877 ( .A(KEYINPUT34), .B(n790), .Z(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U879 ( .A(KEYINPUT36), .B(n793), .ZN(n902) );
  NOR2_X1 U880 ( .A1(n829), .A2(n902), .ZN(n934) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n831) );
  NAND2_X1 U882 ( .A1(n934), .A2(n831), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(KEYINPUT90), .ZN(n827) );
  NAND2_X1 U884 ( .A1(G107), .A2(n895), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(KEYINPUT92), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G95), .A2(n537), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G131), .A2(n889), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G119), .A2(n523), .ZN(n800) );
  XNOR2_X1 U890 ( .A(KEYINPUT91), .B(n800), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT93), .B(n805), .Z(n871) );
  AND2_X1 U894 ( .A1(n871), .A2(G1991), .ZN(n815) );
  XOR2_X1 U895 ( .A(KEYINPUT38), .B(KEYINPUT94), .Z(n807) );
  NAND2_X1 U896 ( .A1(G105), .A2(n537), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n807), .B(n806), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G129), .A2(n523), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G117), .A2(n895), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U901 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n889), .A2(G141), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n872) );
  AND2_X1 U904 ( .A1(n872), .A2(G1996), .ZN(n814) );
  NOR2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n930) );
  INV_X1 U906 ( .A(n831), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n930), .A2(n816), .ZN(n824) );
  INV_X1 U908 ( .A(n824), .ZN(n817) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U910 ( .A1(n984), .A2(n831), .ZN(n818) );
  OR2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n834) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n872), .ZN(n938) );
  NOR2_X1 U913 ( .A1(n871), .A2(G1991), .ZN(n821) );
  XNOR2_X1 U914 ( .A(n821), .B(KEYINPUT104), .ZN(n933) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U916 ( .A1(n933), .A2(n822), .ZN(n823) );
  NOR2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n938), .A2(n825), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT39), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n829), .A2(n902), .ZN(n944) );
  NAND2_X1 U922 ( .A1(n830), .A2(n944), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(n836) );
  XOR2_X1 U925 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n835) );
  XNOR2_X1 U926 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n837), .ZN(G217) );
  NAND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n838) );
  XOR2_X1 U929 ( .A(KEYINPUT106), .B(n838), .Z(n839) );
  NAND2_X1 U930 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U933 ( .A(n842), .ZN(G319) );
  XOR2_X1 U934 ( .A(G1966), .B(G1981), .Z(n844) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U936 ( .A(n844), .B(n843), .ZN(n854) );
  XOR2_X1 U937 ( .A(KEYINPUT111), .B(G2474), .Z(n846) );
  XNOR2_X1 U938 ( .A(G1971), .B(KEYINPUT109), .ZN(n845) );
  XNOR2_X1 U939 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U940 ( .A(G1956), .B(G1961), .Z(n848) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1976), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U943 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U945 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U946 ( .A(n854), .B(n853), .Z(G229) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U948 ( .A(G2072), .B(G2678), .ZN(n855) );
  XNOR2_X1 U949 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U950 ( .A(n857), .B(KEYINPUT42), .Z(n859) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n858) );
  XNOR2_X1 U952 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(G2100), .Z(n861) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U956 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U957 ( .A1(n523), .A2(G124), .ZN(n864) );
  XNOR2_X1 U958 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U959 ( .A1(G112), .A2(n895), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U961 ( .A1(G100), .A2(n537), .ZN(n868) );
  NAND2_X1 U962 ( .A1(G136), .A2(n889), .ZN(n867) );
  NAND2_X1 U963 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U964 ( .A1(n870), .A2(n869), .ZN(G162) );
  XOR2_X1 U965 ( .A(n872), .B(n871), .Z(n873) );
  XNOR2_X1 U966 ( .A(n873), .B(n929), .ZN(n887) );
  XOR2_X1 U967 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U970 ( .A(n876), .B(G162), .Z(n885) );
  NAND2_X1 U971 ( .A1(G103), .A2(n537), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G139), .A2(n889), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U974 ( .A1(G127), .A2(n523), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G115), .A2(n895), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U978 ( .A1(n883), .A2(n882), .ZN(n946) );
  XNOR2_X1 U979 ( .A(G164), .B(n946), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U981 ( .A(n887), .B(n886), .Z(n901) );
  NAND2_X1 U982 ( .A1(n537), .A2(G106), .ZN(n888) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n888), .Z(n891) );
  NAND2_X1 U984 ( .A1(n889), .A2(G142), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n892), .B(KEYINPUT45), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G130), .A2(n523), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U989 ( .A1(n895), .A2(G118), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT112), .B(n896), .Z(n897) );
  NOR2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U992 ( .A(G160), .B(n899), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U994 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U995 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n987), .B(n905), .ZN(n908) );
  XNOR2_X1 U997 ( .A(G171), .B(n906), .ZN(n907) );
  XNOR2_X1 U998 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U999 ( .A(n909), .B(G286), .ZN(n910) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1004 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1007 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1008 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1009 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n919), .ZN(n928) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n928), .ZN(n922) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n924), .A2(n923), .ZN(G225) );
  XOR2_X1 U1017 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1019 ( .A(G120), .ZN(G236) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U1024 ( .A(G261), .ZN(G325) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n928), .ZN(G401) );
  XNOR2_X1 U1027 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1037) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G2090), .B(G162), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n937), .B(KEYINPUT117), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT51), .B(n940), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(KEYINPUT118), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n951) );
  XOR2_X1 U1040 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT50), .B(n949), .Z(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1045 ( .A(KEYINPUT52), .B(n952), .Z(n953) );
  NOR2_X1 U1046 ( .A1(KEYINPUT55), .A2(n953), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT119), .B(n954), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n955), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1049 ( .A(G1991), .B(G25), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n964) );
  XOR2_X1 U1052 ( .A(G2067), .B(G26), .Z(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G28), .ZN(n962) );
  XOR2_X1 U1054 ( .A(KEYINPUT120), .B(n959), .Z(n960) );
  XNOR2_X1 U1055 ( .A(G32), .B(n960), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G27), .B(n965), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1060 ( .A(KEYINPUT53), .B(n968), .Z(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT54), .B(G34), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G2084), .B(n969), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G35), .B(G2090), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(KEYINPUT55), .B(n974), .ZN(n976) );
  INV_X1 U1067 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(G11), .ZN(n1033) );
  XNOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1071 ( .A(G303), .B(G1971), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT125), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G299), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n987), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n1003) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT122), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(n990), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1961), .B(KEYINPUT123), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n992), .B(G301), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT124), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(G168), .B(G1966), .Z(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT121), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n999), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1031) );
  INV_X1 U1093 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1094 ( .A(G1966), .B(G21), .Z(n1013) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G22), .B(G1971), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1099 ( .A(G1986), .B(G24), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1026) );
  XOR2_X1 U1103 ( .A(G1961), .B(G5), .Z(n1024) );
  XNOR2_X1 U1104 ( .A(G20), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G1981), .B(G6), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1015) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(KEYINPUT59), .B(G1348), .Z(n1019) );
  XNOR2_X1 U1110 ( .A(G4), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(n1022), .B(KEYINPUT60), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(n1037), .B(n1036), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

