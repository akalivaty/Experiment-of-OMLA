//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT66), .Z(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G238), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G77), .A2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n213), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n223), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n201), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT68), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  OAI21_X1  g0047(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G150), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n227), .A2(G33), .ZN(new_n251));
  OR2_X1    g0051(.A1(KEYINPUT8), .A2(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT8), .A2(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n248), .B(new_n250), .C1(new_n251), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT70), .B1(new_n210), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n226), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n229), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n260), .A2(new_n264), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n261), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT69), .A2(G223), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT69), .A2(G223), .ZN(new_n273));
  OAI21_X1  g0073(.A(G1698), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n256), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G222), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n284), .C1(G77), .C2(new_n278), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n283), .A2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G226), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G200), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n269), .A2(new_n270), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n271), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT10), .B1(new_n295), .B2(KEYINPUT74), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n269), .B(new_n302), .C1(G179), .C2(new_n292), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G232), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G1698), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(G226), .B2(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(KEYINPUT75), .A3(new_n310), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n284), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n288), .B1(new_n290), .B2(G238), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT76), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  OAI221_X1 g0124(.A(G169), .B1(new_n321), .B2(new_n322), .C1(new_n318), .C2(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G179), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n263), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n334), .A2(new_n262), .A3(G13), .A4(G20), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n331), .B(new_n216), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n249), .A2(G50), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n337), .B1(new_n338), .B2(new_n251), .C1(new_n216), .C2(new_n227), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n260), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n342), .A3(new_n260), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n336), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n260), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(KEYINPUT73), .A3(new_n333), .A4(new_n335), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n333), .A2(new_n335), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n260), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n331), .B1(new_n350), .B2(new_n267), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n332), .B(new_n344), .C1(new_n351), .C2(new_n202), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n330), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(G77), .A3(new_n267), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n338), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n252), .A2(new_n249), .A3(new_n253), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G20), .A2(G77), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n357), .C1(new_n251), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n260), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n362), .A3(new_n260), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n354), .A2(new_n355), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G238), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n278), .B(new_n366), .C1(new_n305), .C2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n284), .C1(G107), .C2(new_n278), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n290), .A2(G244), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n289), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n301), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(G179), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n353), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n370), .A2(new_n293), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(G200), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n365), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n254), .B1(new_n262), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n266), .A2(new_n380), .B1(new_n264), .B2(new_n254), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n249), .A2(G159), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT65), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G68), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(G58), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n205), .A3(new_n203), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n388), .B2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n307), .A2(new_n308), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n227), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR4_X1   g0192(.A1(new_n307), .A2(new_n308), .A3(new_n392), .A4(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n394), .A3(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n260), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n216), .B1(new_n391), .B2(new_n393), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT16), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n381), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G223), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n279), .ZN(new_n401));
  INV_X1    g0201(.A(G226), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(new_n403), .C1(new_n307), .C2(new_n308), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n283), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n283), .A2(G232), .A3(new_n286), .ZN(new_n408));
  NOR4_X1   g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n288), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(new_n405), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n284), .ZN(new_n412));
  INV_X1    g0212(.A(new_n408), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n289), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G169), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n399), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n412), .A2(new_n293), .A3(new_n289), .A4(new_n413), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n406), .A2(new_n288), .A3(new_n408), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(G200), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n381), .C1(new_n396), .C2(new_n398), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n384), .A2(new_n386), .A3(G58), .ZN(new_n429));
  OAI21_X1  g0229(.A(G20), .B1(new_n429), .B2(new_n206), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n382), .ZN(new_n431));
  INV_X1    g0231(.A(new_n216), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n392), .B1(new_n278), .B2(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n428), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n260), .A3(new_n395), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n381), .A4(new_n424), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n421), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n318), .A2(new_n319), .A3(new_n293), .ZN(new_n441));
  INV_X1    g0241(.A(G200), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n327), .B2(new_n328), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n441), .A2(new_n443), .A3(new_n352), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n304), .A2(new_n379), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT83), .ZN(new_n446));
  INV_X1    g0246(.A(G257), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n279), .ZN(new_n448));
  INV_X1    g0248(.A(G264), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G1698), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n450), .C1(new_n307), .C2(new_n308), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT82), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n451), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n284), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT77), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(new_n462), .A3(new_n464), .A4(G274), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n464), .A3(new_n462), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(new_n283), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(G270), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n301), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n283), .ZN(new_n471));
  INV_X1    g0271(.A(G270), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n451), .A2(new_n455), .A3(new_n452), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n455), .B1(new_n451), .B2(new_n452), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(new_n284), .ZN(new_n477));
  AOI22_X1  g0277(.A1(KEYINPUT21), .A2(new_n470), .B1(new_n477), .B2(G179), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n256), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n349), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n348), .A2(new_n260), .A3(new_n347), .ZN(new_n482));
  OAI211_X1 g0282(.A(G116), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  INV_X1    g0286(.A(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n227), .C1(G33), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n260), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n485), .A4(new_n488), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n491), .A2(new_n492), .B1(new_n484), .B2(new_n348), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n483), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n446), .B1(new_n478), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n470), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n498), .B(new_n301), .C1(new_n457), .C2(new_n469), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n457), .A2(new_n469), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n407), .ZN(new_n502));
  OAI211_X1 g0302(.A(KEYINPUT83), .B(new_n494), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(G200), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n477), .A2(G190), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n496), .A2(new_n499), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT84), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n227), .A2(KEYINPUT23), .A3(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT23), .B1(new_n227), .B2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(KEYINPUT23), .C1(new_n227), .C2(G107), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n227), .B(G87), .C1(new_n307), .C2(new_n308), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n509), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n516), .B(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n509), .A4(new_n515), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n260), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n266), .A2(new_n480), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(G107), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n262), .A2(new_n529), .A3(G13), .A4(G20), .ZN(new_n530));
  XOR2_X1   g0330(.A(new_n530), .B(KEYINPUT25), .Z(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G250), .B(new_n279), .C1(new_n307), .C2(new_n308), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n278), .A2(KEYINPUT86), .A3(G250), .A4(new_n279), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G294), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n284), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n468), .A2(G264), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n465), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(new_n284), .B1(G264), .B2(new_n468), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(G190), .A3(new_n465), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n525), .A2(new_n533), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n278), .A2(new_n227), .A3(G68), .ZN(new_n548));
  INV_X1    g0348(.A(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n487), .A3(new_n529), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n310), .A2(new_n227), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT19), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n251), .A2(new_n487), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n552), .C1(KEYINPUT19), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n260), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n348), .A2(new_n358), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n526), .C2(new_n549), .ZN(new_n557));
  INV_X1    g0357(.A(G244), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G1698), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n559), .B1(G238), .B2(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G116), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n283), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n464), .B1(new_n283), .B2(G250), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n262), .A2(G45), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(G274), .ZN(new_n565));
  OR3_X1    g0365(.A1(new_n563), .A2(KEYINPUT80), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT80), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(G190), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n567), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n563), .A2(KEYINPUT80), .A3(new_n565), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n560), .A2(new_n561), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n283), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n543), .A2(new_n301), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n545), .A2(new_n407), .A3(new_n465), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n345), .B1(new_n520), .B2(new_n523), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n532), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n555), .B(new_n556), .C1(new_n358), .C2(new_n526), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(KEYINPUT81), .A3(new_n407), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n573), .B2(new_n301), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n573), .A2(G179), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n580), .B(new_n581), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n547), .A2(new_n575), .A3(new_n579), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n507), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n278), .B2(G250), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n279), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(G1698), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n591), .B(G244), .C1(new_n308), .C2(new_n307), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n558), .B1(new_n276), .B2(new_n277), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n486), .C1(new_n593), .C2(KEYINPUT4), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n284), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n465), .B1(new_n471), .B2(new_n447), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  OAI21_X1  g0399(.A(G244), .B1(new_n307), .B2(new_n308), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n588), .B1(G33), .B2(G283), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n592), .C1(new_n279), .C2(new_n589), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n602), .B2(new_n284), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G190), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n263), .A2(G97), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n529), .A2(KEYINPUT6), .A3(G97), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n487), .A2(new_n529), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(KEYINPUT6), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  OAI21_X1  g0411(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n249), .A2(G77), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n605), .B1(new_n614), .B2(new_n260), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n527), .A2(G97), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n599), .A2(new_n604), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n595), .A2(G179), .A3(new_n597), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n603), .B2(new_n301), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n260), .ZN(new_n620));
  INV_X1    g0420(.A(new_n605), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n616), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT78), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n619), .B2(new_n622), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n622), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT78), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT79), .A3(new_n617), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n445), .A2(new_n587), .A3(new_n628), .A4(new_n633), .ZN(G372));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n570), .B2(new_n571), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n562), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT87), .B1(new_n572), .B2(new_n283), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n636), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n569), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n494), .B1(new_n500), .B2(new_n502), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n499), .A2(new_n579), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n632), .A2(new_n646), .A3(new_n547), .A4(new_n617), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n618), .B(new_n649), .C1(new_n301), .C2(new_n603), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n648), .A2(new_n622), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n644), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n641), .A2(new_n301), .ZN(new_n655));
  INV_X1    g0455(.A(new_n584), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n580), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n575), .A2(new_n630), .A3(new_n585), .A4(new_n631), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n445), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n427), .A2(new_n438), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n374), .A2(new_n661), .A3(new_n444), .ZN(new_n662));
  AOI221_X4 g0462(.A(new_n418), .B1(new_n410), .B2(new_n415), .C1(new_n437), .C2(new_n381), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT18), .B1(new_n399), .B2(new_n416), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n299), .B(new_n300), .C1(new_n662), .C2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n303), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(G369));
  NAND2_X1  g0468(.A1(new_n499), .A2(new_n645), .ZN(new_n669));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n262), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n495), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n669), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n507), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT91), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(KEYINPUT91), .A3(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n678), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n677), .B1(new_n578), .B2(new_n532), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n547), .A2(new_n579), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT92), .B1(new_n579), .B2(new_n678), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n496), .A2(new_n499), .A3(new_n503), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n694), .A3(new_n678), .ZN(new_n695));
  INV_X1    g0495(.A(new_n579), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n678), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  INV_X1    g0500(.A(new_n211), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(G41), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n211), .A2(KEYINPUT93), .A3(new_n461), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n550), .A2(G116), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n262), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n230), .B2(new_n705), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND2_X1  g0509(.A1(new_n647), .A2(new_n653), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n643), .ZN(new_n711));
  INV_X1    g0511(.A(new_n659), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n677), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n587), .A2(new_n628), .A3(new_n633), .A4(new_n678), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n641), .A2(new_n407), .A3(new_n501), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n543), .A2(new_n719), .A3(new_n598), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n543), .B2(new_n598), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n477), .A2(G179), .A3(new_n545), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n603), .A2(new_n568), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n598), .A2(new_n573), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n502), .A3(KEYINPUT30), .A4(new_n545), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n677), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n677), .C1(new_n722), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n716), .B1(new_n717), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n617), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n630), .B2(new_n631), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n496), .A2(new_n579), .A3(new_n499), .A4(new_n503), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n547), .A4(new_n643), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n624), .A2(new_n625), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(new_n652), .A3(new_n575), .A4(new_n585), .ZN(new_n742));
  INV_X1    g0542(.A(new_n657), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n643), .A2(new_n622), .A3(new_n648), .A4(new_n650), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(KEYINPUT26), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n678), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT29), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n715), .A2(new_n736), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n709), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n687), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n262), .B1(new_n671), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n705), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n752), .B(new_n756), .C1(G330), .C2(new_n682), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n227), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n407), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n758), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n390), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n442), .A2(G179), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(G20), .A2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n765), .B1(new_n771), .B2(G303), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(new_n769), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G322), .ZN(new_n775));
  NAND3_X1  g0575(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n293), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G326), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n227), .B1(new_n759), .B2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(G294), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n767), .A2(new_n758), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G283), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n772), .A2(new_n775), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n764), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G77), .B1(G50), .B2(new_n777), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n201), .B2(new_n773), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT96), .ZN(new_n793));
  INV_X1    g0593(.A(new_n760), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n783), .A2(new_n487), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n793), .B(new_n798), .C1(new_n549), .C2(new_n770), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n278), .B1(new_n202), .B2(new_n780), .C1(new_n786), .C2(new_n529), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n789), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n226), .B1(G20), .B2(new_n301), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n230), .A2(new_n463), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n390), .A2(new_n211), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(new_n243), .C2(new_n463), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n278), .A2(G355), .A3(new_n211), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G116), .C2(new_n211), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n802), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n756), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n812), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n803), .B(new_n814), .C1(new_n682), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n757), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n373), .A2(KEYINPUT100), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT100), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n365), .A2(new_n820), .A3(new_n372), .A4(new_n371), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n377), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n678), .B(new_n822), .C1(new_n654), .C2(new_n659), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n373), .A2(new_n678), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n365), .A2(new_n677), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n823), .B1(new_n713), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(new_n736), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n736), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n756), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n802), .A2(new_n810), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n755), .B1(G77), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT98), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n774), .A2(G143), .B1(G150), .B2(new_n779), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(new_n777), .ZN(new_n838));
  INV_X1    g0638(.A(G159), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n836), .B1(new_n837), .B2(new_n838), .C1(new_n839), .C2(new_n764), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n278), .B1(new_n843), .B2(new_n760), .C1(new_n770), .C2(new_n229), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n840), .A2(new_n841), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n787), .A2(G68), .B1(G58), .B2(new_n784), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n764), .A2(new_n484), .ZN(new_n849));
  INV_X1    g0649(.A(G303), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n838), .A2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n797), .B(new_n851), .C1(G283), .C2(new_n779), .ZN(new_n852));
  INV_X1    g0652(.A(G294), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n390), .B1(new_n760), .B2(new_n762), .C1(new_n853), .C2(new_n773), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n787), .B2(G87), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n852), .B(new_n855), .C1(new_n529), .C2(new_n770), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n848), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n835), .B1(new_n857), .B2(new_n802), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT99), .ZN(new_n859));
  INV_X1    g0659(.A(new_n826), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n811), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n831), .A2(new_n861), .ZN(G384));
  AOI21_X1  g0662(.A(new_n409), .B1(G169), .B2(new_n414), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n437), .A2(new_n381), .B1(new_n863), .B2(new_n675), .ZN(new_n864));
  INV_X1    g0664(.A(new_n425), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT104), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n675), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n399), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT104), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n417), .A2(new_n868), .A3(new_n869), .A4(new_n425), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n868), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n665), .B2(new_n661), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n866), .A2(new_n870), .A3(new_n874), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT16), .B1(new_n389), .B2(new_n394), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n381), .B1(new_n396), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n867), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n665), .B2(new_n661), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n872), .B1(new_n864), .B2(new_n865), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n416), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT37), .A4(new_n425), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n717), .A2(new_n734), .ZN(new_n894));
  INV_X1    g0694(.A(new_n444), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n352), .A2(new_n677), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n353), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n352), .B(new_n677), .C1(new_n330), .C2(new_n444), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n826), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n894), .A4(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n885), .B1(new_n421), .B2(new_n439), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n888), .A2(new_n890), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n881), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n892), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n894), .A3(new_n907), .A4(new_n899), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT105), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n901), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n445), .A2(new_n894), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G330), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n906), .A2(new_n907), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT39), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n893), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n353), .A2(new_n677), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n897), .A2(new_n898), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n819), .A2(new_n678), .A3(new_n821), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n823), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n907), .A3(new_n906), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n665), .A2(new_n675), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n715), .A2(new_n748), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n445), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n667), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n931), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n918), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n262), .B2(new_n671), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n484), .B1(new_n610), .B2(KEYINPUT35), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n228), .C1(KEYINPUT35), .C2(new_n610), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n230), .A2(G77), .A3(new_n387), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(G50), .B2(new_n202), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n670), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(new_n940), .A3(new_n943), .ZN(G367));
  NAND2_X1  g0744(.A1(new_n622), .A2(new_n677), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n738), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n651), .A2(new_n677), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n695), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT42), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n741), .B1(new_n948), .B2(new_n696), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n678), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n557), .A2(new_n677), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n657), .A2(new_n643), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n657), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n961), .A2(new_n687), .A3(new_n692), .A4(new_n948), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n956), .C1(new_n693), .C2(new_n949), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n704), .B(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n698), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT45), .B1(new_n698), .B2(new_n948), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT44), .B1(new_n698), .B2(new_n948), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n948), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n693), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n973), .C1(new_n970), .C2(new_n971), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n687), .A3(new_n692), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n694), .A2(new_n678), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n692), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n687), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n685), .A2(new_n686), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n975), .A2(new_n977), .A3(new_n750), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n969), .B1(new_n984), .B2(new_n750), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n965), .B(new_n967), .C1(new_n985), .C2(new_n754), .ZN(new_n986));
  INV_X1    g0786(.A(G150), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n278), .B1(new_n760), .B2(new_n837), .C1(new_n987), .C2(new_n773), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n771), .B2(G58), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n790), .A2(G50), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n777), .A2(G143), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n780), .B2(new_n839), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G68), .B2(new_n784), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n787), .A2(G77), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n771), .A2(G116), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n390), .B1(new_n760), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n786), .A2(new_n487), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G283), .C2(new_n790), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n838), .A2(new_n762), .B1(new_n783), .B2(new_n529), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G294), .B2(new_n779), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n773), .A2(new_n850), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT109), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n756), .B1(new_n1008), .B2(new_n802), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n806), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n813), .B1(new_n211), .B2(new_n358), .C1(new_n1010), .C2(new_n238), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(new_n815), .C2(new_n959), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT110), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n986), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n750), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n981), .A2(new_n749), .A3(new_n982), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n705), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n774), .A2(G317), .B1(G311), .B2(new_n779), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n777), .A2(G322), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n850), .C2(new_n764), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1021), .B1(new_n1022), .B2(new_n783), .C1(new_n853), .C2(new_n770), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n794), .A2(G326), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n278), .B1(new_n787), .B2(G116), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n390), .B1(new_n790), .B2(G68), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n229), .B2(new_n773), .C1(new_n987), .C2(new_n760), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n770), .A2(new_n338), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n783), .A2(new_n358), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n838), .B2(new_n839), .C1(new_n254), .C2(new_n780), .ZN(new_n1034));
  OR4_X1    g0834(.A1(new_n1000), .A2(new_n1031), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n756), .B1(new_n1036), .B2(new_n802), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n254), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n229), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n706), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n463), .C1(KEYINPUT50), .C2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G68), .B2(G77), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n806), .B1(new_n235), .B2(new_n463), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n706), .A2(new_n211), .A3(new_n278), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n211), .A2(G107), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n813), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n692), .A2(new_n815), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1037), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n983), .B2(new_n754), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1017), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1017), .A2(KEYINPUT111), .A3(new_n1050), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n975), .A2(new_n977), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n1015), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n705), .A3(new_n984), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n975), .A2(new_n754), .A3(new_n977), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G87), .A2(new_n787), .B1(new_n771), .B2(new_n216), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n794), .A2(G143), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n838), .A2(new_n987), .B1(new_n773), .B2(new_n839), .ZN(new_n1062));
  XOR2_X1   g0862(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n783), .A2(new_n338), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n278), .B1(new_n764), .B2(new_n254), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n779), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n780), .A2(new_n850), .B1(new_n783), .B2(new_n484), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n278), .B(new_n1069), .C1(G322), .C2(new_n794), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G107), .A2(new_n787), .B1(new_n771), .B2(G283), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n853), .C2(new_n764), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n838), .A2(new_n998), .B1(new_n773), .B2(new_n762), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1068), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n802), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n806), .A2(new_n246), .B1(G97), .B2(new_n701), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n813), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n755), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT114), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n815), .B2(new_n948), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1058), .A2(new_n1059), .A3(new_n1082), .ZN(G390));
  AOI21_X1  g0883(.A(new_n921), .B1(new_n906), .B2(new_n907), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT39), .B1(new_n882), .B2(new_n892), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n928), .A2(new_n923), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n746), .A2(new_n678), .A3(new_n822), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n927), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n925), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n923), .B1(new_n882), .B2(new_n892), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n735), .A2(new_n899), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT115), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1086), .A2(new_n1094), .A3(new_n1091), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n754), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n810), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n786), .A2(new_n202), .B1(new_n853), .B2(new_n760), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT118), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n390), .B1(new_n770), .B2(new_n549), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n774), .A2(G116), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n780), .A2(new_n529), .B1(new_n838), .B2(new_n1022), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1065), .B(new_n1106), .C1(G97), .C2(new_n790), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT119), .Z(new_n1109));
  NOR2_X1   g0909(.A1(new_n773), .A2(new_n843), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n770), .A2(new_n987), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n780), .A2(new_n837), .B1(new_n838), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G159), .B2(new_n784), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n278), .B1(new_n760), .B2(new_n1116), .C1(new_n764), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n787), .B2(G50), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1112), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1109), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n756), .B1(new_n1121), .B2(new_n802), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1100), .B(new_n1122), .C1(new_n1038), .C2(new_n833), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1099), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n925), .B1(new_n827), .B2(new_n735), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1125), .A2(new_n1093), .A3(new_n1088), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n735), .A2(new_n860), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n926), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n735), .A2(new_n899), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1127), .A2(KEYINPUT116), .A3(new_n926), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n823), .A2(new_n927), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1126), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n933), .B(new_n667), .C1(new_n716), .C2(new_n916), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n704), .B1(new_n1137), .B2(new_n1098), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1136), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n1131), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT116), .B1(new_n1127), .B2(new_n926), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1126), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1086), .A2(new_n1094), .A3(new_n1091), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1094), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1124), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G378));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n304), .B(KEYINPUT120), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n269), .A2(new_n867), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n1157), .A3(new_n1152), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G330), .B(new_n900), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n931), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n914), .B2(G330), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1164), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n931), .A2(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n911), .A2(new_n913), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1173), .A3(G330), .A4(new_n900), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1174), .A3(new_n1163), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n754), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n794), .A2(G283), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n529), .B2(new_n773), .C1(new_n358), .C2(new_n764), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n786), .A2(new_n201), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n390), .A2(new_n461), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1179), .A2(new_n1032), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n784), .A2(G68), .B1(G116), .B2(new_n777), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n487), .C2(new_n780), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT58), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n229), .B1(new_n307), .B2(G41), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n780), .A2(new_n843), .B1(new_n783), .B2(new_n987), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n838), .A2(new_n1116), .B1(new_n773), .B2(new_n1113), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n837), .B2(new_n764), .C1(new_n770), .C2(new_n1117), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT59), .Z(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(new_n787), .B2(G159), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G33), .B1(new_n794), .B2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1185), .A2(new_n1186), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n756), .B1(new_n1195), .B2(new_n802), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(G50), .B2(new_n833), .C1(new_n1164), .C2(new_n811), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1177), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1139), .B1(new_n1148), .B2(new_n1135), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1172), .A2(new_n1174), .A3(new_n1163), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1163), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1201));
  OAI211_X1 g1001(.A(KEYINPUT57), .B(new_n1199), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT121), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1176), .A2(new_n1204), .A3(KEYINPUT57), .A4(new_n1199), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1136), .B1(new_n1098), .B2(new_n1144), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n705), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1198), .B1(new_n1206), .B2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n969), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1145), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n201), .A2(new_n786), .B1(new_n770), .B2(new_n839), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n278), .B1(new_n783), .B2(new_n229), .C1(new_n987), .C2(new_n764), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n777), .A2(G132), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G137), .A2(new_n774), .B1(new_n1216), .B2(KEYINPUT122), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(KEYINPUT122), .B2(new_n1216), .C1(new_n780), .C2(new_n1117), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1214), .B(new_n1215), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .C1(new_n1113), .C2(new_n760), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n760), .A2(new_n850), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1033), .B1(new_n838), .B2(new_n853), .C1(new_n484), .C2(new_n780), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n390), .B1(new_n773), .B2(new_n1022), .C1(new_n529), .C2(new_n764), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n787), .B2(G77), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(new_n487), .C2(new_n770), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1221), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n756), .B1(new_n1228), .B2(new_n802), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n925), .B2(new_n811), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n202), .B2(new_n832), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1144), .B2(new_n754), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(G381));
  NAND3_X1  g1033(.A1(new_n1150), .A2(new_n1177), .A3(new_n1197), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n704), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1053), .A2(new_n817), .A3(new_n1054), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(G387), .A2(new_n1241), .A3(G390), .A4(G381), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  NAND4_X1  g1046(.A1(new_n1136), .A2(new_n1142), .A3(new_n1143), .A4(KEYINPUT60), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1145), .A2(new_n1247), .A3(new_n705), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT60), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1232), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1243), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G384), .B(new_n1232), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n676), .A2(G213), .A3(G2897), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1254), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1150), .B1(new_n1239), .B2(new_n1198), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n676), .A2(G213), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1234), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1259), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1251), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1257), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(new_n1256), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT63), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1260), .A2(new_n1264), .A3(new_n1253), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1274), .A2(KEYINPUT125), .A3(new_n1241), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n986), .A2(G390), .A3(new_n1013), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G390), .B1(new_n986), .B2(new_n1013), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1241), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1277), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1279), .B(new_n1280), .C1(new_n1283), .C2(new_n1275), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(KEYINPUT63), .B2(new_n1271), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1273), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1271), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1280), .B1(new_n1289), .B2(new_n1268), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1260), .A2(new_n1264), .A3(KEYINPUT62), .A4(new_n1253), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1279), .B1(new_n1283), .B2(new_n1275), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1286), .B1(new_n1292), .B2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(G378), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1245), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1240), .B2(new_n1260), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1253), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT126), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1293), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1301), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1240), .A2(new_n1260), .A3(KEYINPUT127), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1297), .B1(new_n1296), .B2(new_n1245), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1294), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1304), .A2(new_n1310), .ZN(G402));
endmodule


