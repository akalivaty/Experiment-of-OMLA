//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G122), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G122), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n189), .B(new_n191), .C1(KEYINPUT14), .C2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n190), .B2(G122), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n190), .A2(G122), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n188), .A2(G116), .ZN(new_n196));
  OAI211_X1 g010(.A(G107), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT67), .A2(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(G143), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT65), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT65), .A2(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n202), .B2(new_n207), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n193), .B(new_n197), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n211));
  INV_X1    g025(.A(new_n201), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT67), .A2(G128), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT13), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n199), .B2(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(KEYINPUT13), .A3(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G134), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n189), .A2(new_n191), .A3(G107), .ZN(new_n221));
  AOI21_X1  g035(.A(G107), .B1(new_n189), .B2(new_n191), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n210), .A2(new_n211), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n211), .B1(new_n210), .B2(new_n225), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT9), .B(G234), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G217), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n197), .A2(new_n193), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT65), .A2(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT65), .A2(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n215), .B2(new_n206), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n235), .B1(new_n224), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT92), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n210), .A2(new_n211), .A3(new_n225), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n233), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n232), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT93), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n231), .B1(new_n226), .B2(new_n227), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n233), .A3(new_n242), .ZN(new_n248));
  AOI21_X1  g062(.A(G902), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT93), .ZN(new_n250));
  INV_X1    g064(.A(G478), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(KEYINPUT15), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n252), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT94), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n246), .A2(new_n250), .A3(KEYINPUT94), .A4(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(G214), .B1(G237), .B2(G902), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G210), .B1(G237), .B2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  INV_X1    g077(.A(G113), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n190), .A2(G119), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G119), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G116), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n190), .A2(G119), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT5), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(KEYINPUT2), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G113), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G116), .B(G119), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G104), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(new_n280), .B2(G107), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n192), .A3(G104), .ZN(new_n283));
  INV_X1    g097(.A(G101), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(G107), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(new_n283), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n280), .A2(G107), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n192), .A2(G104), .ZN(new_n288));
  OAI21_X1  g102(.A(G101), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n286), .A2(KEYINPUT4), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n281), .A2(new_n283), .A3(new_n285), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G101), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n276), .B1(new_n277), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n269), .A2(new_n270), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n273), .A4(new_n275), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n292), .A2(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n300), .A3(G101), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n293), .A2(new_n303), .A3(new_n300), .A4(G101), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n291), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G110), .B(G122), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n263), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n291), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n302), .A2(new_n304), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n286), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n298), .A2(new_n296), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n307), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT0), .A2(G128), .ZN(new_n319));
  XNOR2_X1  g133(.A(G143), .B(G146), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(KEYINPUT64), .ZN(new_n321));
  INV_X1    g135(.A(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G143), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n214), .A2(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT0), .A2(G128), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT64), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n318), .B1(new_n330), .B2(G125), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n200), .A2(new_n201), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n323), .A2(new_n324), .A3(G128), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n336), .A2(new_n325), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n318), .A3(new_n341), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT85), .Z(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n320), .B1(new_n334), .B2(new_n335), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n323), .A2(new_n324), .A3(G128), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n338), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT84), .A4(G125), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n342), .B2(new_n331), .ZN(new_n354));
  INV_X1    g168(.A(new_n348), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n314), .A2(new_n263), .A3(new_n315), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n317), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n286), .A2(new_n289), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(KEYINPUT87), .A3(new_n278), .A4(new_n272), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n307), .B(KEYINPUT8), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n361), .A2(KEYINPUT87), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n286), .A2(new_n289), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n279), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n343), .A2(new_n344), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n307), .B(new_n309), .C1(new_n310), .C2(new_n313), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(KEYINPUT89), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT7), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n347), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n373), .B(new_n374), .C1(new_n354), .C2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n187), .B1(new_n370), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n262), .B1(new_n359), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n368), .B(KEYINPUT88), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n345), .A2(new_n375), .A3(new_n378), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n374), .A3(new_n373), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n317), .A2(new_n357), .A3(new_n358), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n187), .A4(new_n261), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n260), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n280), .ZN(new_n390));
  INV_X1    g204(.A(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n341), .A2(G140), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n341), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n394), .A2(G146), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(G146), .B1(new_n394), .B2(new_n395), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G237), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n230), .A3(G214), .ZN(new_n400));
  NOR2_X1   g214(.A1(KEYINPUT90), .A2(G143), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(G237), .A2(G953), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(G214), .C1(KEYINPUT90), .C2(G143), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT17), .A3(G131), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n398), .B(new_n406), .C1(new_n410), .C2(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(KEYINPUT18), .A3(G131), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n392), .A2(new_n393), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(G146), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT18), .A2(G131), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n402), .A2(new_n404), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n390), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n409), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n408), .B1(new_n402), .B2(new_n404), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n394), .A2(new_n395), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n322), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n394), .A2(new_n395), .A3(G146), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n406), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n390), .B(new_n417), .C1(new_n421), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n411), .A2(KEYINPUT91), .A3(new_n390), .A4(new_n417), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n418), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G475), .B1(new_n430), .B2(G902), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n230), .A2(G952), .ZN(new_n432));
  INV_X1    g246(.A(G234), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n399), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n187), .B(new_n230), .C1(G234), .C2(G237), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(G898), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n429), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n413), .B(KEYINPUT19), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n410), .B(new_n424), .C1(G146), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n417), .ZN(new_n444));
  INV_X1    g258(.A(new_n390), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(G475), .A2(G902), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n428), .A2(new_n429), .B1(new_n445), .B2(new_n444), .ZN(new_n450));
  INV_X1    g264(.A(new_n448), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n431), .B(new_n439), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n258), .A2(new_n388), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G140), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n230), .A2(G227), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT11), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G137), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n460), .A2(new_n203), .A3(new_n204), .ZN(new_n461));
  INV_X1    g275(.A(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT11), .A3(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n461), .A2(G131), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(KEYINPUT11), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n236), .A2(new_n468), .A3(new_n237), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n408), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n311), .A2(new_n321), .A3(new_n329), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n310), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n330), .B1(new_n294), .B2(new_n292), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n305), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n337), .A2(new_n339), .ZN(new_n478));
  INV_X1    g292(.A(new_n324), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n325), .A2(new_n199), .B1(new_n479), .B2(KEYINPUT1), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n290), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT10), .B1(new_n350), .B2(new_n352), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n481), .A2(KEYINPUT10), .B1(new_n482), .B2(new_n290), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n471), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n471), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n486), .B(new_n483), .C1(new_n474), .C2(new_n476), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n458), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT83), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n305), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT80), .B1(new_n475), .B2(new_n305), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n471), .B(new_n484), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n458), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n290), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n497), .A2(new_n350), .A3(new_n352), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n486), .B1(new_n498), .B2(new_n481), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT12), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(KEYINPUT82), .A3(new_n493), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n504), .B(new_n458), .C1(new_n485), .C2(new_n487), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G469), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n187), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n458), .B1(new_n500), .B2(new_n487), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n477), .A2(new_n484), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n486), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n494), .B2(KEYINPUT81), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n492), .B2(new_n493), .ZN(new_n514));
  OAI211_X1 g328(.A(G469), .B(new_n509), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(G469), .A2(G902), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G221), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n229), .B2(new_n187), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n520), .B(KEYINPUT78), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n455), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n321), .B(new_n329), .C1(new_n466), .C2(new_n470), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n469), .A2(new_n408), .A3(new_n463), .A4(new_n464), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n408), .B1(G134), .B2(G137), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n238), .B2(G137), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(new_n527), .C1(new_n350), .C2(new_n352), .ZN(new_n528));
  INV_X1    g342(.A(new_n312), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n470), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n330), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n527), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n340), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT30), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n536), .A3(new_n528), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n530), .B1(new_n538), .B2(new_n312), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n403), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT29), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n529), .B1(new_n524), .B2(new_n528), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT28), .B1(new_n530), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT69), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT70), .B1(new_n532), .B2(new_n534), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n524), .A2(new_n551), .A3(new_n528), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n529), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n548), .A2(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n530), .C2(new_n547), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n544), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n546), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n530), .B2(new_n547), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n554), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n544), .A2(KEYINPUT29), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n559), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND4_X1   g383(.A1(new_n559), .A2(new_n565), .A3(new_n566), .A4(new_n568), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n558), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G472), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  INV_X1    g387(.A(new_n537), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n536), .B1(new_n524), .B2(new_n528), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n312), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n530), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n544), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n539), .A2(new_n580), .A3(new_n544), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT71), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n548), .A2(new_n549), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n556), .A3(new_n566), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n545), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n579), .A4(new_n581), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n573), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT32), .B(new_n593), .C1(new_n584), .C2(new_n589), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n572), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G217), .B1(new_n433), .B2(G902), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT74), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n424), .B1(G146), .B2(new_n413), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT24), .B(G110), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n212), .A2(new_n213), .A3(new_n268), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n199), .A2(G119), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n602), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .A4(new_n201), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT75), .ZN(new_n607));
  INV_X1    g421(.A(G110), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT75), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n599), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  INV_X1    g428(.A(new_n602), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n335), .B2(new_n268), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n600), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n398), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT76), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n599), .ZN(new_n620));
  INV_X1    g434(.A(new_n612), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n603), .A2(new_n609), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n614), .ZN(new_n624));
  OAI221_X1 g438(.A(new_n624), .B1(new_n616), .B2(new_n600), .C1(new_n396), .C2(new_n397), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT76), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT22), .B(G137), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n519), .A2(new_n433), .A3(G953), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n619), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n623), .A2(new_n625), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT76), .A3(new_n630), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT25), .B1(new_n635), .B2(new_n187), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT25), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n637), .B(G902), .C1(new_n632), .C2(new_n634), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n598), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n596), .A2(new_n187), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT77), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n523), .A2(new_n595), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  AOI21_X1  g459(.A(new_n593), .B1(new_n584), .B2(new_n589), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n590), .A2(new_n187), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(G472), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n521), .B1(new_n508), .B2(new_n517), .ZN(new_n649));
  INV_X1    g463(.A(new_n388), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n438), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n648), .A2(new_n643), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n451), .B1(new_n441), .B2(new_n446), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n440), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT20), .B1(new_n450), .B2(new_n451), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n431), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n247), .A2(new_n248), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n247), .A2(KEYINPUT33), .A3(new_n248), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(G478), .A3(new_n187), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n652), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  INV_X1    g482(.A(new_n258), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n655), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g485(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n450), .C2(new_n451), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n653), .B2(new_n440), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n450), .A2(KEYINPUT96), .A3(KEYINPUT20), .A4(new_n451), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n671), .B(new_n672), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n431), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(KEYINPUT97), .B(G475), .C1(new_n430), .C2(G902), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n651), .A2(new_n669), .A3(new_n676), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(new_n643), .A3(new_n649), .A4(new_n648), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT35), .B(G107), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n632), .A2(new_n634), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n637), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n635), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n597), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n631), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n633), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n641), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n686), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n639), .A2(KEYINPUT98), .A3(new_n693), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n523), .A2(new_n648), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  INV_X1    g514(.A(new_n436), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n434), .B1(new_n701), .B2(G900), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT99), .Z(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n678), .A2(new_n679), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n676), .A3(new_n256), .A4(new_n257), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT100), .B1(new_n706), .B2(new_n650), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n705), .A2(new_n676), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n388), .A4(new_n669), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n595), .A3(new_n649), .A4(new_n697), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT101), .B(G128), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G30));
  XOR2_X1   g528(.A(new_n703), .B(KEYINPUT39), .Z(new_n715));
  NAND2_X1  g529(.A1(new_n649), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n187), .B1(new_n564), .B2(new_n544), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n539), .A2(new_n545), .ZN(new_n720));
  OAI21_X1  g534(.A(G472), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n592), .B2(new_n594), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n382), .A2(new_n387), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT38), .Z(new_n724));
  AND2_X1   g538(.A1(new_n656), .A2(new_n431), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n258), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n259), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n724), .A2(new_n727), .A3(new_n697), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n717), .A2(new_n718), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  AOI22_X1  g544(.A1(new_n656), .A2(new_n431), .B1(new_n658), .B2(new_n663), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n704), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n650), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n595), .A2(new_n649), .A3(new_n697), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NAND2_X1  g549(.A1(new_n506), .A2(new_n187), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  INV_X1    g551(.A(new_n520), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n508), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n737), .A2(KEYINPUT102), .A3(new_n738), .A4(new_n508), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n595), .A3(new_n643), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n651), .A2(new_n731), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT41), .B(G113), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NOR2_X1   g561(.A1(new_n743), .A2(new_n681), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n190), .ZN(G18));
  NAND3_X1  g563(.A1(new_n741), .A2(new_n388), .A3(new_n742), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n669), .A2(new_n453), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n595), .A2(new_n751), .A3(new_n697), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n268), .ZN(G21));
  AOI21_X1  g568(.A(new_n580), .B1(new_n539), .B2(new_n544), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n529), .B1(new_n535), .B2(new_n537), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n545), .A4(new_n530), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n567), .B2(new_n544), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n591), .B(KEYINPUT103), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(G902), .B1(new_n584), .B2(new_n589), .ZN(new_n762));
  INV_X1    g576(.A(G472), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n643), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n726), .A2(new_n388), .A3(new_n439), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n741), .A3(new_n742), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT104), .B(G122), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G24));
  AND3_X1   g583(.A1(new_n506), .A2(new_n507), .A3(new_n187), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n507), .B1(new_n506), .B2(new_n187), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT102), .B1(new_n772), .B2(new_n738), .ZN(new_n773));
  INV_X1    g587(.A(new_n742), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n639), .A2(KEYINPUT98), .A3(new_n693), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT98), .B1(new_n639), .B2(new_n693), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n647), .A2(G472), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT105), .A3(new_n697), .A4(new_n761), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n704), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT106), .B1(new_n731), .B2(new_n704), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n784), .A3(new_n388), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G125), .ZN(G27));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n595), .A2(new_n643), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n382), .A2(new_n259), .A3(new_n387), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n520), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n518), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n787), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n790), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n794), .A2(new_n786), .A3(new_n785), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT42), .A3(new_n643), .A4(new_n595), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  OR2_X1    g615(.A1(new_n794), .A2(new_n706), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n791), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(G134), .Z(G36));
  NAND2_X1  g618(.A1(new_n725), .A2(new_n664), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT43), .Z(new_n806));
  NOR3_X1   g620(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT71), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n588), .B1(new_n758), .B2(new_n587), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n591), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n782), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT107), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n697), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n811), .B1(new_n810), .B2(new_n697), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT45), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n507), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n516), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n508), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n738), .B(new_n715), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n792), .B(KEYINPUT108), .Z(new_n829));
  NAND2_X1  g643(.A1(new_n815), .A2(new_n816), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n817), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  OAI21_X1  g646(.A(new_n738), .B1(new_n825), .B2(new_n826), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(KEYINPUT109), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(KEYINPUT109), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n595), .A2(new_n643), .A3(new_n732), .A4(new_n792), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n837), .B(new_n838), .C1(new_n833), .C2(new_n836), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G140), .ZN(G42));
  AND2_X1   g654(.A1(new_n781), .A2(new_n783), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n741), .A2(new_n388), .A3(new_n787), .A4(new_n742), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n650), .A2(new_n258), .A3(new_n725), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n703), .B(KEYINPUT114), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n690), .A2(new_n520), .A3(new_n694), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n722), .A2(new_n518), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n712), .A2(new_n734), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT115), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n649), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n809), .A2(KEYINPUT32), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n646), .A2(new_n573), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n853), .B2(new_n572), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n854), .B(new_n697), .C1(new_n711), .C2(new_n733), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n788), .A2(new_n855), .A3(new_n856), .A4(new_n847), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n743), .A2(new_n681), .B1(new_n750), .B2(new_n752), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n767), .B1(new_n743), .B2(new_n744), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n803), .B1(new_n797), .B2(new_n799), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n256), .A2(KEYINPUT110), .A3(new_n257), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT110), .B1(new_n256), .B2(new_n257), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n863), .B(new_n725), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n665), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT110), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT94), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n244), .B2(new_n252), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT93), .B1(new_n659), .B2(new_n187), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n245), .B(G902), .C1(new_n247), .C2(new_n248), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n873), .B2(new_n252), .ZN(new_n874));
  INV_X1    g688(.A(new_n257), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n256), .A2(KEYINPUT110), .A3(new_n257), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n863), .B1(new_n878), .B2(new_n725), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n644), .B(new_n698), .C1(new_n880), .C2(new_n652), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n796), .B1(new_n781), .B2(new_n783), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n885));
  INV_X1    g699(.A(new_n792), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n708), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n887), .B2(new_n878), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n705), .A2(new_n676), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n792), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT112), .A3(new_n877), .A4(new_n876), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n595), .A2(new_n649), .A3(new_n697), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n888), .A2(new_n891), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n854), .A2(new_n895), .A3(KEYINPUT113), .A4(new_n697), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n861), .A2(new_n862), .A3(new_n883), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n858), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n849), .A2(new_n857), .A3(KEYINPUT52), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(new_n848), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n788), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n858), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n905), .B2(KEYINPUT53), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n858), .A2(new_n898), .A3(new_n911), .A4(new_n904), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT53), .B1(new_n899), .B2(new_n900), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n849), .A2(new_n857), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n902), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n861), .A2(new_n862), .A3(new_n883), .A4(new_n897), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n900), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n919), .B2(new_n911), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n909), .B(new_n910), .C1(KEYINPUT54), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n806), .A2(new_n435), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n764), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n260), .A2(new_n925), .A3(new_n724), .A4(new_n775), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n928));
  NOR4_X1   g742(.A1(new_n773), .A2(new_n774), .A3(new_n434), .A4(new_n792), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n806), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n927), .A2(new_n928), .B1(new_n784), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n837), .B1(new_n833), .B2(new_n836), .ZN(new_n932));
  INV_X1    g746(.A(new_n772), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n522), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n829), .A3(new_n925), .ZN(new_n935));
  INV_X1    g749(.A(new_n722), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n643), .A3(new_n936), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n937), .A2(new_n657), .A3(new_n664), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT51), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n925), .A2(new_n388), .A3(new_n775), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(new_n432), .C1(new_n937), .C2(new_n665), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT118), .ZN(new_n945));
  INV_X1    g759(.A(new_n791), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n930), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT48), .Z(new_n948));
  NOR2_X1   g762(.A1(new_n944), .A2(KEYINPUT118), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n941), .A2(new_n942), .A3(new_n945), .A4(new_n950), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n923), .A2(new_n951), .B1(G952), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n772), .B(KEYINPUT49), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n805), .A2(new_n521), .A3(new_n260), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n724), .A2(new_n954), .A3(new_n643), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n936), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(G75));
  NOR2_X1   g771(.A1(new_n230), .A2(G952), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n922), .A2(G210), .A3(G902), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n317), .A2(new_n358), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n357), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT55), .Z(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT119), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n962), .A2(new_n969), .A3(new_n965), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(G51));
  XOR2_X1   g785(.A(new_n516), .B(KEYINPUT57), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n919), .A2(new_n914), .A3(new_n911), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n905), .A2(KEYINPUT53), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n975), .A2(KEYINPUT54), .A3(new_n920), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT54), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n915), .B2(new_n921), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n972), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT120), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(KEYINPUT120), .B(new_n972), .C1(new_n976), .C2(new_n978), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n506), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n975), .A2(new_n920), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n984), .A2(new_n187), .A3(new_n821), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n958), .B1(new_n983), .B2(new_n985), .ZN(G54));
  NAND4_X1  g800(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n450), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n450), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n958), .ZN(G60));
  AND2_X1   g804(.A1(new_n661), .A2(new_n662), .ZN(new_n991));
  NAND2_X1  g805(.A1(G478), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT59), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n923), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n976), .A2(new_n978), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n991), .A2(new_n993), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n959), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n994), .A2(new_n997), .ZN(G63));
  NAND2_X1  g812(.A1(G217), .A2(G902), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT121), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT60), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n922), .A2(new_n692), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n922), .A2(new_n1001), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n959), .B(new_n1002), .C1(new_n1003), .C2(new_n635), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G66));
  NOR3_X1   g820(.A1(new_n859), .A2(new_n860), .A3(new_n881), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(G953), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT122), .ZN(new_n1009));
  OAI21_X1  g823(.A(G953), .B1(new_n437), .B2(new_n346), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n963), .B1(G898), .B2(new_n230), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(G69));
  AND2_X1   g827(.A1(new_n831), .A2(new_n839), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n828), .A2(new_n946), .A3(new_n844), .ZN(new_n1015));
  INV_X1    g829(.A(new_n862), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n788), .A2(new_n855), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(G953), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n230), .A2(G900), .ZN(new_n1020));
  OAI21_X1  g834(.A(KEYINPUT123), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT123), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1020), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1018), .A2(new_n831), .A3(new_n839), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(G953), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n538), .B(new_n442), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1021), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  OR4_X1    g842(.A1(new_n791), .A2(new_n880), .A3(new_n716), .A4(new_n792), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n831), .A2(new_n839), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n788), .A2(new_n729), .A3(new_n855), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT62), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n230), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT124), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n230), .B1(G227), .B2(G900), .ZN(new_n1035));
  AOI22_X1  g849(.A1(new_n1033), .A2(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT125), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1035), .A2(new_n1034), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT125), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1028), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1039), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(G72));
  INV_X1    g858(.A(new_n720), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  NOR2_X1   g861(.A1(new_n540), .A2(new_n544), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n906), .A2(new_n1045), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1047), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1051), .B1(new_n1024), .B2(new_n1007), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1050), .B(new_n959), .C1(new_n1052), .C2(new_n1049), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n1007), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n1047), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(KEYINPUT126), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT126), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1055), .A2(new_n1058), .A3(new_n1047), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1057), .A2(new_n720), .A3(new_n1059), .ZN(new_n1060));
  OR2_X1    g874(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1053), .B1(new_n1061), .B2(new_n1062), .ZN(G57));
endmodule


