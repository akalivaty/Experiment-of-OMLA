//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G97), .B(G107), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G41), .A2(G45), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT65), .B1(new_n254), .B2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT65), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n256), .B(new_n208), .C1(G41), .C2(G45), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G222), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n263), .B1(new_n264), .B2(new_n261), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(new_n218), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT66), .B1(new_n271), .B2(new_n251), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n260), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(KEYINPUT68), .B(G179), .Z(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n218), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(KEYINPUT67), .A2(KEYINPUT8), .A3(G58), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT8), .B1(KEYINPUT67), .B2(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n209), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n278), .B1(new_n208), .B2(G20), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G50), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n276), .B(new_n296), .C1(G169), .C2(new_n274), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n295), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(KEYINPUT70), .A3(KEYINPUT9), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n274), .A2(G190), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n274), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n303), .B2(new_n302), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n306), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n297), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT7), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n261), .A2(new_n315), .A3(G20), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n209), .ZN(new_n322));
  OAI21_X1  g0122(.A(G68), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n222), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n325), .B2(new_n201), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n286), .A2(G159), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(KEYINPUT16), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n315), .B1(new_n261), .B2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n222), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n334), .B2(new_n328), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n278), .ZN(new_n336));
  INV_X1    g0136(.A(new_n294), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n282), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n290), .A2(new_n209), .A3(G1), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n282), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n255), .A2(G232), .A3(new_n252), .A4(new_n257), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n253), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n318), .A2(new_n320), .A3(G226), .A4(G1698), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n318), .A2(new_n320), .A3(G223), .A4(new_n262), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n347), .B(new_n348), .C1(new_n317), .C2(new_n224), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n273), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n275), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n350), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n342), .A2(new_n344), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT18), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n342), .A2(new_n357), .A3(new_n344), .A4(new_n354), .ZN(new_n358));
  INV_X1    g0158(.A(new_n346), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n349), .A2(new_n273), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n350), .B2(G200), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(new_n336), .A3(new_n340), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n363), .A2(new_n336), .A3(KEYINPUT17), .A4(new_n340), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n356), .A2(new_n358), .A3(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT12), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n339), .B2(new_n222), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n370), .A2(new_n372), .B1(new_n337), .B2(new_n222), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n264), .B2(new_n283), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT11), .B1(new_n375), .B2(new_n278), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  INV_X1    g0182(.A(new_n258), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n250), .A2(new_n252), .A3(new_n385), .A4(G274), .ZN(new_n386));
  AOI22_X1  g0186(.A1(G238), .A2(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n318), .A2(new_n320), .A3(G232), .A4(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n318), .A2(new_n320), .A3(G226), .A4(new_n262), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n273), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n382), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n384), .A2(new_n386), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n255), .A2(G238), .A3(new_n252), .A4(new_n257), .ZN(new_n395));
  AND4_X1   g0195(.A1(new_n382), .A2(new_n392), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n381), .B(G169), .C1(new_n393), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n387), .A2(new_n382), .A3(new_n392), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(G179), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n381), .B1(new_n403), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n380), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(G200), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n379), .C1(new_n361), .C2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G107), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n265), .A2(new_n223), .B1(new_n409), .B2(new_n261), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n261), .A2(G232), .A3(new_n262), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n273), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n252), .A2(G274), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n383), .A2(G244), .B1(new_n250), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G200), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n339), .A2(new_n264), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n337), .B2(new_n264), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT8), .B(G58), .Z(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n284), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n279), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n416), .B(new_n425), .C1(new_n361), .C2(new_n415), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n415), .A2(new_n353), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n412), .A2(new_n275), .A3(new_n414), .ZN(new_n428));
  INV_X1    g0228(.A(new_n425), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NOR4_X1   g0231(.A1(new_n314), .A2(new_n369), .A3(new_n408), .A4(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT23), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n409), .A3(G20), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT78), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n433), .A2(new_n435), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n318), .A2(new_n320), .A3(new_n209), .A4(G87), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT22), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT22), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n261), .A2(new_n444), .A3(new_n209), .A4(G87), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT24), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n441), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n441), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n278), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n249), .A2(G1), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n252), .ZN(new_n455));
  INV_X1    g0255(.A(G264), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT79), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n451), .B1(new_n271), .B2(new_n251), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT79), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(G264), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n318), .A2(new_n320), .A3(G257), .A4(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n318), .A2(new_n320), .A3(G250), .A4(new_n262), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G294), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n457), .A2(new_n461), .B1(new_n273), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n208), .A2(G45), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n413), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(G190), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n273), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n459), .B2(G264), .ZN(new_n474));
  AND4_X1   g0274(.A1(new_n460), .A2(new_n454), .A3(G264), .A4(new_n252), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n208), .A2(G33), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n279), .A2(new_n292), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n409), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT25), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n292), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n339), .A2(KEYINPUT25), .A3(new_n409), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND4_X1   g0284(.A1(new_n450), .A2(new_n472), .A3(new_n477), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n476), .A2(G169), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  INV_X1    g0289(.A(G179), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n476), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n466), .A2(KEYINPUT81), .A3(G179), .A4(new_n471), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n476), .A2(KEYINPUT80), .A3(G169), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n488), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n450), .A2(new_n484), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n277), .A2(new_n218), .B1(G20), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n209), .C1(G33), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT76), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT76), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n498), .A2(new_n505), .A3(new_n501), .A4(KEYINPUT20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n479), .A2(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n292), .A2(new_n497), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n318), .A2(new_n320), .A3(G264), .A4(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n318), .A2(new_n320), .A3(G257), .A4(new_n262), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n261), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n273), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n459), .A2(G270), .B1(new_n413), .B2(new_n470), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n353), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n518), .A3(G190), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n508), .A3(new_n511), .A4(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(new_n518), .A3(G179), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n512), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n512), .A2(new_n519), .A3(new_n530), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n522), .A2(new_n526), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(new_n262), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n499), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G250), .A2(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT4), .A2(G244), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n261), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n273), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n252), .A2(new_n269), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n271), .A2(KEYINPUT66), .A3(new_n251), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n535), .B2(new_n540), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n454), .A2(G257), .A3(new_n252), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n471), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n543), .A2(new_n549), .A3(new_n275), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n471), .A2(new_n550), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n353), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n286), .A2(G77), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n556), .A2(new_n500), .A3(G107), .ZN(new_n557));
  XNOR2_X1  g0357(.A(G97), .B(G107), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(new_n559), .B2(new_n209), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n409), .B1(new_n332), .B2(new_n333), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n278), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  MUX2_X1   g0362(.A(new_n292), .B(new_n479), .S(G97), .Z(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n552), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n541), .A2(new_n548), .A3(new_n273), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n548), .B1(new_n541), .B2(new_n273), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n308), .B1(new_n568), .B2(new_n551), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n547), .A2(new_n553), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n562), .A3(new_n563), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n565), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(G1698), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n318), .A2(new_n320), .A3(G238), .A4(new_n262), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G116), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n273), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n451), .A2(new_n225), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n413), .A2(new_n451), .B1(new_n252), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(new_n580), .A3(new_n275), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n578), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT75), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n224), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G97), .A2(G107), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT74), .A2(G87), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n209), .B1(new_n390), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n318), .A2(new_n320), .A3(new_n209), .A4(G68), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n283), .B2(new_n500), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n278), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n421), .A2(new_n339), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n479), .A2(new_n421), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n584), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n595), .A2(new_n278), .B1(new_n339), .B2(new_n421), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n584), .B1(new_n600), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n583), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n479), .A2(new_n224), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n578), .A2(new_n580), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n579), .A2(new_n252), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n252), .A2(G274), .A3(new_n451), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n577), .B2(new_n273), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G190), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n573), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n432), .A2(new_n496), .A3(new_n532), .A4(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n297), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n341), .A2(new_n354), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT18), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n341), .A2(new_n354), .A3(new_n357), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n430), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n407), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n405), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n366), .A2(new_n367), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n312), .A2(new_n313), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n617), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n432), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n522), .A2(new_n529), .A3(new_n531), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n495), .B2(new_n494), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n596), .A2(new_n598), .A3(new_n597), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT75), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n600), .A2(new_n584), .A3(new_n598), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n606), .A2(new_n361), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n604), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n636), .A2(new_n583), .B1(new_n638), .B2(new_n607), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n450), .A2(new_n472), .A3(new_n477), .A4(new_n484), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n543), .A2(new_n549), .A3(new_n551), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  INV_X1    g0442(.A(new_n564), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(new_n571), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n639), .A2(new_n640), .A3(new_n565), .A4(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n602), .B1(new_n632), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n614), .A2(new_n647), .A3(new_n565), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT82), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n471), .A2(new_n550), .A3(new_n275), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n566), .A2(new_n567), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n554), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n552), .A2(KEYINPUT82), .A3(new_n554), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n564), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(KEYINPUT83), .B(new_n647), .C1(new_n655), .C2(new_n614), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n647), .B1(new_n655), .B2(new_n614), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT83), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n646), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n629), .B1(new_n630), .B2(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n291), .A2(new_n209), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(G213), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n512), .A2(new_n668), .ZN(new_n669));
  MUX2_X1   g0469(.A(new_n532), .B(new_n631), .S(new_n669), .Z(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n495), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n496), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n494), .A2(new_n495), .A3(new_n668), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n522), .A2(new_n529), .A3(new_n531), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n668), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n496), .ZN(new_n684));
  INV_X1    g0484(.A(new_n668), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n494), .A2(new_n495), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT84), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n681), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n212), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n589), .A2(G116), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n216), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g0496(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n661), .B2(new_n668), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n552), .A2(new_n554), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n643), .B1(new_n701), .B2(new_n649), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n639), .A2(new_n702), .A3(KEYINPUT26), .A4(new_n654), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n647), .B1(new_n614), .B2(new_n565), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n685), .B1(new_n646), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT88), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  INV_X1    g0507(.A(new_n602), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n573), .A2(new_n614), .A3(new_n485), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n494), .A2(new_n495), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n682), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n703), .A2(new_n704), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n668), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n700), .A2(new_n707), .A3(new_n716), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n496), .A2(new_n615), .A3(new_n532), .A4(new_n685), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n466), .A2(new_n570), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n528), .A4(new_n611), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n351), .B1(new_n517), .B2(new_n518), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n641), .A2(new_n476), .A3(new_n606), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n466), .A2(new_n570), .A3(new_n611), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n527), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n668), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n528), .A2(new_n466), .A3(new_n570), .A4(new_n611), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n721), .A2(new_n476), .A3(new_n606), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n723), .A2(new_n730), .B1(new_n731), .B2(new_n641), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n685), .B1(new_n732), .B2(new_n720), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n733), .B2(KEYINPUT31), .ZN(new_n734));
  OAI21_X1  g0534(.A(G330), .B1(new_n718), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n717), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n698), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n290), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT89), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n249), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n693), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT90), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT90), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n673), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n671), .A2(new_n672), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n671), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n690), .A2(new_n321), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G355), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G116), .B2(new_n212), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n243), .A2(new_n249), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n690), .A2(new_n261), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n249), .B2(new_n217), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n754), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n218), .B1(G20), .B2(new_n353), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT92), .Z(new_n763));
  OAI21_X1  g0563(.A(new_n745), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT95), .B1(new_n490), .B2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n209), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n490), .A2(KEYINPUT95), .A3(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G20), .A3(new_n490), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT94), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n261), .B1(new_n779), .B2(G329), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n768), .A2(new_n361), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n515), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n275), .A2(new_n209), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n772), .B(new_n783), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT93), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n784), .A2(new_n789), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n773), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n361), .A2(G200), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n791), .B2(new_n792), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n794), .B1(new_n797), .B2(G322), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n785), .A2(new_n361), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n209), .B1(new_n795), .B2(new_n490), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G326), .B1(G294), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n788), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n586), .A2(new_n588), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n781), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n779), .A2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(new_n786), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(KEYINPUT32), .C1(new_n808), .C2(new_n222), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n324), .A2(new_n796), .B1(new_n793), .B2(new_n264), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n807), .A2(KEYINPUT32), .ZN(new_n811));
  INV_X1    g0611(.A(new_n799), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n202), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n261), .B1(new_n500), .B2(new_n800), .C1(new_n770), .C2(new_n409), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n804), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n764), .B1(new_n816), .B2(new_n761), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n746), .A2(new_n747), .B1(new_n751), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n430), .A2(KEYINPUT102), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n429), .A2(new_n668), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT102), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n427), .A2(new_n429), .A3(new_n822), .A4(new_n428), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n426), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n623), .A2(new_n668), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n661), .B2(new_n668), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n648), .A2(new_n656), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n639), .A2(new_n702), .A3(new_n654), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT83), .B1(new_n830), .B2(new_n647), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n712), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n820), .A2(new_n426), .A3(new_n823), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n685), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n744), .B1(new_n837), .B2(new_n735), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n735), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(KEYINPUT103), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT103), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n779), .A2(G132), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n769), .A2(G68), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n781), .A2(G50), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n321), .B1(new_n801), .B2(G58), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G137), .A2(new_n799), .B1(new_n786), .B2(G150), .ZN(new_n847));
  INV_X1    g0647(.A(G159), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT99), .B(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n793), .C1(new_n796), .C2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT100), .Z(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n771), .A2(new_n808), .B1(new_n812), .B2(new_n515), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n794), .B2(G116), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT97), .Z(new_n857));
  NAND2_X1  g0657(.A1(new_n769), .A2(G87), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n778), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT98), .Z(new_n861));
  OAI221_X1 g0661(.A(new_n321), .B1(new_n500), .B2(new_n800), .C1(new_n782), .C2(new_n409), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n797), .B2(G294), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n857), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  INV_X1    g0666(.A(new_n761), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n761), .A2(new_n748), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n745), .B1(G77), .B2(new_n870), .C1(new_n826), .C2(new_n749), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n841), .B1(new_n868), .B2(new_n871), .ZN(G384));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n615), .A2(new_n496), .A3(new_n532), .A4(new_n685), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n728), .B1(new_n726), .B2(new_n668), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n380), .A2(new_n668), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n408), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n879), .B(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n405), .A3(new_n407), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n878), .A2(new_n885), .A3(new_n826), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(new_n666), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n342), .A2(new_n344), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n355), .A2(new_n889), .A3(new_n890), .A4(new_n364), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n364), .A2(KEYINPUT106), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n363), .A2(new_n336), .A3(new_n894), .A4(new_n340), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n618), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT107), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT107), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n893), .A2(new_n898), .A3(new_n618), .A4(new_n895), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n892), .B1(new_n900), .B2(KEYINPUT37), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT108), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n621), .B1(new_n902), .B2(new_n368), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n626), .A2(KEYINPUT108), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n889), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n887), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n666), .B1(new_n336), .B2(new_n340), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n618), .A2(new_n364), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n908), .B2(new_n907), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n369), .A2(new_n907), .B1(new_n909), .B2(new_n891), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT38), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n873), .B(new_n886), .C1(new_n906), .C2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n878), .A2(new_n885), .A3(new_n826), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n369), .A2(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n891), .A2(new_n909), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n873), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n432), .A2(new_n878), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n672), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n405), .A2(new_n668), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT39), .B1(new_n917), .B2(new_n916), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n899), .A2(new_n889), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n364), .A2(KEYINPUT106), .B1(new_n341), .B2(new_n354), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n898), .B1(new_n929), .B2(new_n895), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT37), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n366), .A2(new_n902), .A3(new_n367), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n622), .A2(new_n904), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n889), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n931), .A2(new_n891), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n911), .B(new_n927), .C1(new_n935), .C2(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n925), .B1(new_n926), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n660), .A2(new_n648), .A3(new_n656), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n834), .B1(new_n938), .B2(new_n712), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n820), .A2(new_n823), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n685), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT104), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n885), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n917), .A2(new_n916), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n944), .A2(new_n945), .B1(new_n622), .B2(new_n888), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n700), .A2(new_n707), .A3(new_n432), .A4(new_n716), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n629), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n924), .A2(new_n950), .B1(G1), .B2(new_n739), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n924), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(new_n559), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(G116), .A3(new_n219), .A4(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n216), .A2(new_n264), .A3(new_n325), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n222), .A2(G50), .ZN(new_n959));
  OAI211_X1 g0759(.A(G1), .B(new_n290), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT110), .ZN(G367));
  NAND3_X1  g0762(.A1(new_n702), .A2(new_n654), .A3(new_n668), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n644), .B(new_n565), .C1(new_n643), .C2(new_n685), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n565), .B1(new_n966), .B2(new_n710), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n685), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n684), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT42), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT112), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n605), .A2(new_n685), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n708), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n614), .B2(new_n972), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n971), .B(new_n974), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n968), .A2(new_n970), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT43), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n681), .B2(new_n966), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n681), .A2(new_n966), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(KEYINPUT43), .C2(new_n975), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n691), .B(KEYINPUT41), .Z(new_n982));
  INV_X1    g0782(.A(new_n965), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n688), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT45), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n687), .A2(KEYINPUT84), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n983), .B1(KEYINPUT113), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n687), .A2(KEYINPUT84), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(KEYINPUT113), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n680), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n678), .A2(new_n683), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT114), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n684), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n673), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n736), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n982), .B1(new_n1003), .B2(new_n736), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n740), .A2(new_n208), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n979), .B(new_n981), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n757), .A2(new_n239), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n763), .B1(new_n690), .B2(new_n422), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n744), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n750), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n769), .A2(G97), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n261), .B1(new_n801), .B2(G107), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n1013), .C1(new_n1014), .C2(new_n778), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n782), .A2(new_n497), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n771), .B2(new_n793), .ZN(new_n1018));
  INV_X1    g0818(.A(G294), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n808), .B1(new_n812), .B2(new_n859), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n796), .A2(new_n515), .B1(new_n1016), .B2(KEYINPUT46), .ZN(new_n1021));
  OR4_X1    g0821(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n770), .A2(new_n264), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n808), .B2(new_n848), .C1(new_n812), .C2(new_n849), .ZN(new_n1025));
  INV_X1    g0825(.A(G137), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n261), .B1(new_n222), .B2(new_n800), .C1(new_n778), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G58), .B2(new_n781), .ZN(new_n1028));
  INV_X1    g0828(.A(G150), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n202), .B2(new_n793), .C1(new_n1029), .C2(new_n796), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1022), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1010), .B1(new_n1011), .B2(new_n974), .C1(new_n1032), .C2(new_n867), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1007), .A2(new_n1033), .ZN(G387));
  AOI22_X1  g0834(.A1(G311), .A2(new_n786), .B1(new_n799), .B2(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n515), .B2(new_n793), .C1(new_n1014), .C2(new_n796), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n781), .A2(G294), .B1(G283), .B2(new_n801), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT49), .Z(new_n1042));
  AOI21_X1  g0842(.A(new_n261), .B1(new_n779), .B2(G326), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n497), .B2(new_n770), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n812), .A2(new_n848), .B1(new_n264), .B2(new_n782), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n779), .A2(G150), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n801), .A2(new_n422), .ZN(new_n1048));
  AND4_X1   g0848(.A1(new_n261), .A2(new_n1047), .A3(new_n1012), .A4(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n202), .B2(new_n796), .C1(new_n222), .C2(new_n793), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1046), .B(new_n1050), .C1(new_n282), .C2(new_n786), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n761), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n419), .A2(new_n202), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT50), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n758), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n249), .B2(new_n236), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n752), .A2(new_n694), .B1(new_n409), .B2(new_n690), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT115), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1052), .B(new_n745), .C1(new_n763), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n679), .B2(new_n750), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1001), .A2(new_n691), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1000), .A2(new_n736), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(G393));
  AOI21_X1  g0866(.A(new_n692), .B1(new_n994), .B2(new_n1002), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1002), .B2(new_n994), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n966), .A2(new_n750), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n758), .A2(new_n246), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n763), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n500), .B2(new_n212), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n745), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n321), .B1(new_n801), .B2(G77), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n858), .B(new_n1074), .C1(new_n778), .C2(new_n849), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n808), .A2(new_n202), .B1(new_n222), .B2(new_n782), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n794), .C2(new_n419), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n796), .A2(new_n848), .B1(new_n812), .B2(new_n1029), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n796), .A2(new_n859), .B1(new_n812), .B2(new_n1014), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n786), .A2(G303), .B1(G116), .B2(new_n801), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n1019), .C2(new_n793), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n261), .B1(new_n779), .B2(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n409), .B2(new_n770), .C1(new_n771), .C2(new_n782), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT116), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n1080), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1073), .B1(new_n1088), .B2(new_n761), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT117), .Z(new_n1090));
  AOI22_X1  g0890(.A1(new_n994), .A2(new_n1006), .B1(new_n1069), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1068), .A2(new_n1091), .ZN(G390));
  INV_X1    g0892(.A(new_n885), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n943), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n836), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n925), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n926), .B(new_n936), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n685), .B(new_n833), .C1(new_n646), .C2(new_n705), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n885), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n911), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1101), .A3(new_n925), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n827), .B1(new_n881), .B2(new_n884), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n735), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1097), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n876), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n672), .B1(new_n1109), .B2(new_n874), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1103), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n885), .B1(new_n1110), .B2(new_n826), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1105), .A2(new_n1114), .A3(new_n1099), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n826), .C1(new_n718), .C2(new_n734), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1093), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1111), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1094), .B1(new_n661), .B2(new_n834), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1116), .A2(new_n1093), .B1(new_n1110), .B2(new_n1103), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n943), .B1(new_n832), .B2(new_n835), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1115), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n432), .A2(new_n1110), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n948), .A2(new_n629), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n692), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n926), .A2(new_n936), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1096), .B1(new_n1120), .B2(new_n885), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1102), .B(new_n1106), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n907), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n626), .B1(KEYINPUT18), .B2(new_n355), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n358), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n891), .A2(new_n909), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n887), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n911), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT39), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1138), .A2(KEYINPUT39), .B1(new_n906), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n944), .A2(new_n925), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1096), .B1(new_n1099), .B2(new_n885), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1140), .A2(new_n1141), .B1(new_n1101), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1132), .B1(new_n1143), .B2(new_n1111), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n1105), .A2(new_n1114), .A3(new_n1099), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1119), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1122), .A2(KEYINPUT118), .A3(new_n1123), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1127), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT119), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1144), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1129), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1113), .A2(new_n1006), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n745), .B1(new_n282), .B2(new_n870), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n808), .A2(new_n409), .B1(new_n224), .B2(new_n782), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G283), .B2(new_n799), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n794), .A2(G97), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n797), .A2(G116), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n779), .A2(G294), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n261), .B1(new_n801), .B2(G77), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1161), .A2(new_n843), .A3(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n781), .A2(G150), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT120), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT53), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n261), .B1(new_n848), .B2(new_n800), .C1(new_n778), .C2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G50), .B2(new_n769), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n799), .B1(new_n786), .B2(G137), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G132), .A2(new_n797), .B1(new_n794), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .A4(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1166), .A2(KEYINPUT53), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1164), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1156), .B1(new_n1177), .B2(new_n761), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1130), .B2(new_n749), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1155), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1154), .A2(new_n1180), .ZN(G378));
  AOI21_X1  g0981(.A(new_n744), .B1(new_n202), .B2(new_n869), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n793), .A2(new_n1026), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n786), .A2(G132), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n799), .A2(G125), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n801), .A2(G150), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n781), .A2(new_n1173), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1183), .B(new_n1188), .C1(G128), .C2(new_n797), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n769), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n770), .A2(new_n324), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n808), .A2(new_n500), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G116), .C2(new_n799), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n321), .A2(new_n248), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n801), .B2(G68), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n771), .B2(new_n778), .C1(new_n782), .C2(new_n264), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n794), .B2(new_n422), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1198), .B(new_n1202), .C1(new_n409), .C2(new_n796), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1199), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1195), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1209));
  NAND2_X1  g1009(.A1(new_n314), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n302), .A2(new_n888), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  INV_X1    g1012(.A(new_n1209), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n297), .B(new_n1213), .C1(new_n312), .C2(new_n313), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1210), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1212), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1182), .B1(new_n867), .B2(new_n1208), .C1(new_n1217), .C2(new_n749), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT123), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n886), .B1(new_n1137), .B2(new_n911), .ZN(new_n1221));
  OAI21_X1  g1021(.A(G330), .B1(new_n1221), .B2(KEYINPUT40), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n1222), .B2(new_n912), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n672), .B1(new_n918), .B2(new_n873), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1101), .A2(KEYINPUT40), .A3(new_n913), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1217), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n937), .A2(new_n946), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1223), .B2(new_n1227), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1220), .B1(new_n1231), .B2(new_n1006), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1127), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1222), .A2(new_n912), .A3(new_n1217), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1226), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n947), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(KEYINPUT57), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n691), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1149), .B1(new_n1144), .B2(new_n1125), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1232), .B1(new_n1239), .B2(new_n1241), .ZN(G375));
  XNOR2_X1  g1042(.A(new_n1005), .B(KEYINPUT124), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n885), .A2(new_n749), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n808), .A2(new_n497), .B1(new_n500), .B2(new_n782), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G294), .B2(new_n799), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n794), .A2(G107), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n797), .A2(G283), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n321), .B(new_n1048), .C1(new_n778), .C2(new_n515), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1023), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n261), .B1(new_n800), .B2(new_n202), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1252), .B(new_n1196), .C1(G128), .C2(new_n779), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n1026), .B2(new_n796), .C1(new_n1029), .C2(new_n793), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n799), .A2(G132), .B1(G159), .B2(new_n781), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n808), .B2(new_n1172), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1251), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n761), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1258), .B(new_n745), .C1(G68), .C2(new_n870), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1125), .A2(new_n1243), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1128), .A2(new_n982), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(G381));
  OR4_X1    g1064(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1265), .A2(G387), .A3(G381), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1219), .B1(new_n1267), .B2(new_n1005), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1231), .A2(new_n1240), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT57), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1229), .A2(new_n1230), .A3(new_n1270), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n692), .B1(new_n1272), .B2(new_n1240), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1268), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n691), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1107), .A2(new_n1112), .B1(new_n1127), .B2(new_n1125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT119), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1144), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1155), .A2(new_n1179), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1154), .B2(new_n1180), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1266), .A2(new_n1274), .A3(new_n1284), .ZN(G407));
  INV_X1    g1085(.A(G213), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(G343), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1274), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(G213), .A3(new_n1288), .ZN(G409));
  XNOR2_X1  g1089(.A(G393), .B(G396), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G390), .B1(new_n1007), .B2(new_n1033), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1007), .A2(new_n1033), .A3(G390), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(new_n1292), .A3(new_n1290), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(G375), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1302), .A2(KEYINPUT126), .A3(G378), .A4(new_n1232), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  OAI221_X1 g1104(.A(new_n1219), .B1(new_n1267), .B2(new_n1243), .C1(new_n1269), .C2(new_n982), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1284), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1287), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1150), .A2(KEYINPUT60), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1308), .A2(new_n1263), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n692), .B1(new_n1308), .B2(new_n1263), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1260), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(G384), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT62), .B1(new_n1307), .B2(new_n1313), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1301), .A2(new_n1303), .B1(new_n1284), .B2(new_n1305), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NOR4_X1   g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1287), .A4(new_n1312), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1314), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT126), .B1(new_n1274), .B2(G378), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(G375), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1306), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1287), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1313), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(new_n1318), .A3(new_n1316), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1311), .A2(G384), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1311), .A2(G384), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1287), .A2(G2897), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1325), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1298), .B1(new_n1319), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1307), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1324), .A2(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .A4(new_n1333), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(new_n1304), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1274), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1343));
  OR3_X1    g1143(.A1(new_n1342), .A2(new_n1313), .A3(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1313), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1298), .B(new_n1346), .ZN(G402));
endmodule


