//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(new_n458), .A3(KEYINPUT3), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n458), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n459), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n458), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n471), .A2(G136), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n469), .A2(G2105), .A3(new_n462), .A4(new_n460), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n469), .A2(new_n460), .A3(new_n462), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n495));
  NOR4_X1   g070(.A1(new_n474), .A2(KEYINPUT4), .A3(new_n490), .A4(G2105), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n464), .A2(KEYINPUT68), .A3(G114), .ZN(new_n502));
  OAI221_X1 g077(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n509));
  INV_X1    g084(.A(new_n496), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n504), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n505), .A2(new_n513), .ZN(G164));
  XOR2_X1   g089(.A(KEYINPUT6), .B(G651), .Z(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT71), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(G50), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT73), .Z(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(G62), .B2(new_n518), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n521), .A2(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT75), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT76), .B(G51), .Z(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n516), .B(KEYINPUT5), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n515), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G89), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n538), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G651), .B1(new_n540), .B2(G90), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n532), .A2(G543), .A3(new_n534), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n553), .B2(G52), .ZN(G171));
  NAND2_X1  g129(.A1(new_n553), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n539), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n540), .B2(G81), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n535), .A2(KEYINPUT78), .A3(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n539), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n540), .B2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n535), .A2(G49), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n518), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n540), .B2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n539), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(G48), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n539), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(new_n533), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n539), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n540), .B2(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n536), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n553), .A2(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(new_n540), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n539), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n600), .A2(new_n601), .B1(G651), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  XNOR2_X1  g184(.A(G284), .B(KEYINPUT80), .ZN(G321));
  NAND2_X1  g185(.A1(G299), .A2(new_n607), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n471), .A2(G135), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n464), .A2(KEYINPUT82), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT82), .B1(new_n464), .B2(G111), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  AND4_X1   g201(.A1(G2104), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n484), .B2(G123), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n475), .A2(new_n478), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n644), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  INV_X1    g235(.A(new_n657), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n661), .B2(new_n655), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n655), .B(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n662), .B1(new_n664), .B2(new_n661), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n661), .A3(new_n658), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n660), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT20), .Z(new_n679));
  OR2_X1    g254(.A1(new_n672), .A2(new_n674), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(new_n677), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n677), .A3(new_n675), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(G23), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n577), .A2(new_n579), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  MUX2_X1   g277(.A(G6), .B(G305), .S(G16), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n695), .A2(new_n701), .A3(new_n702), .A4(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n484), .A2(G119), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n464), .A2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n471), .A2(KEYINPUT87), .A3(G131), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT87), .B1(new_n471), .B2(G131), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n709), .B1(new_n710), .B2(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G25), .B(new_n714), .S(G29), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT88), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n715), .B(new_n717), .Z(new_n718));
  MUX2_X1   g293(.A(G24), .B(G290), .S(G16), .Z(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1986), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n708), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(KEYINPUT36), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(KEYINPUT36), .C2(new_n724), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n691), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n560), .B2(new_n691), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  NOR2_X1   g309(.A1(G171), .A2(new_n691), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G5), .B2(new_n691), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n739), .B2(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT24), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n480), .B2(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n691), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT23), .Z(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n691), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n614), .B2(new_n691), .ZN(new_n750));
  INV_X1    g325(.A(G1348), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n734), .A2(new_n744), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n691), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n691), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n742), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND4_X1  g334(.A1(new_n463), .A2(G140), .A3(new_n464), .A4(new_n469), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n483), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n759), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n757), .B(new_n769), .C1(new_n737), .C2(new_n736), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n742), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n471), .A2(G139), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(new_n464), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n772), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(new_n742), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G2072), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n484), .A2(G129), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT26), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n784), .A2(new_n785), .B1(G105), .B2(new_n478), .ZN(new_n786));
  INV_X1    g361(.A(G141), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n786), .C1(new_n470), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G29), .B2(G32), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n780), .B(new_n793), .C1(new_n738), .C2(new_n743), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n753), .B(new_n770), .C1(new_n794), .C2(KEYINPUT95), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(KEYINPUT95), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g371(.A1(G164), .A2(new_n742), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G27), .B2(new_n742), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT31), .B(G11), .Z(new_n801));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n742), .B1(new_n802), .B2(G28), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n804), .A2(KEYINPUT96), .B1(new_n802), .B2(G28), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n630), .B2(new_n742), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT97), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n742), .A2(G35), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT98), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G162), .B2(new_n742), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2090), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n809), .B(new_n816), .C1(new_n792), .C2(new_n791), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  INV_X1    g394(.A(new_n798), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(G2078), .B2(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n796), .A2(new_n800), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n730), .A2(new_n731), .A3(new_n822), .ZN(G311));
  NAND3_X1  g398(.A1(new_n730), .A2(new_n731), .A3(new_n822), .ZN(G150));
  NOR2_X1   g399(.A1(new_n606), .A2(new_n615), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n540), .A2(G93), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n526), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n553), .B2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n560), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n555), .A2(new_n559), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n553), .A2(G55), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n830), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n827), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  AOI21_X1  g413(.A(G860), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT102), .Z(new_n841));
  OAI21_X1  g416(.A(G860), .B1(new_n834), .B2(new_n830), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n488), .B(new_n480), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n629), .B(new_n845), .Z(new_n846));
  INV_X1    g421(.A(new_n777), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n511), .A2(new_n512), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n767), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n496), .B1(new_n507), .B2(KEYINPUT69), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n504), .B1(new_n850), .B2(new_n509), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n765), .A2(new_n851), .A3(new_n766), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n788), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  INV_X1    g432(.A(new_n852), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n851), .B1(new_n765), .B2(new_n766), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n789), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n788), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n849), .A2(new_n862), .A3(new_n852), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n857), .B1(new_n864), .B2(new_n778), .ZN(new_n865));
  INV_X1    g440(.A(new_n778), .ZN(new_n866));
  AOI211_X1 g441(.A(KEYINPUT103), .B(new_n866), .C1(new_n860), .C2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n856), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n471), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n484), .A2(G130), .ZN(new_n870));
  OR2_X1    g445(.A1(G106), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n873), .B(new_n856), .C1(new_n865), .C2(new_n867), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n714), .B(new_n634), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n846), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n846), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g462(.A(G288), .B(G303), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G305), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT42), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n614), .A2(new_n567), .A3(new_n571), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(new_n606), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n898), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n836), .B(new_n617), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n902), .B(new_n903), .S(new_n904), .Z(new_n905));
  AOI21_X1  g480(.A(new_n895), .B1(new_n905), .B2(KEYINPUT105), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(KEYINPUT105), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G868), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n831), .ZN(G295));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n831), .ZN(G331));
  NAND3_X1  g486(.A1(new_n832), .A2(G301), .A3(new_n835), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G301), .B1(new_n832), .B2(new_n835), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(G286), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n836), .A2(G171), .ZN(new_n916));
  AOI21_X1  g491(.A(G168), .B1(new_n916), .B2(new_n912), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n903), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(G286), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(G168), .A3(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n902), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n921), .A3(new_n890), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n885), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n901), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT106), .A4(new_n900), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n898), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n898), .B2(KEYINPUT41), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n919), .A2(new_n920), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n918), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n890), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(KEYINPUT43), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n919), .A2(new_n902), .A3(new_n920), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n898), .B1(new_n919), .B2(new_n920), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n885), .A3(new_n922), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n924), .A2(new_n941), .A3(new_n935), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n943), .B1(KEYINPUT44), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n851), .B2(G1384), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(G40), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n472), .A2(new_n477), .A3(new_n479), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G2067), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n767), .B(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n854), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n789), .B2(new_n956), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n714), .B(new_n717), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(G290), .B(G1986), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n953), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT123), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n967));
  INV_X1    g542(.A(new_n952), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT109), .B1(new_n851), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n970), .B(new_n971), .C1(new_n497), .C2(new_n504), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n848), .A2(KEYINPUT70), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n851), .A2(new_n506), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n968), .B(new_n974), .C1(new_n977), .C2(new_n973), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n967), .B1(new_n978), .B2(G2084), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n974), .A2(new_n968), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(KEYINPUT116), .A3(new_n738), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n969), .A2(new_n972), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n952), .B1(new_n984), .B2(new_n948), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT45), .B(new_n971), .C1(new_n505), .C2(new_n513), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n983), .B(G1966), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n970), .B1(new_n848), .B2(new_n971), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT109), .B(G1384), .C1(new_n511), .C2(new_n512), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n948), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n968), .A3(new_n986), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT115), .B1(new_n991), .B2(new_n756), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n979), .B(new_n982), .C1(new_n987), .C2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n964), .B(new_n966), .C1(new_n993), .C2(G286), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(G8), .A3(G286), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n756), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n983), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(KEYINPUT115), .A3(new_n756), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(G168), .A3(new_n979), .A4(new_n982), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n964), .B1(new_n1001), .B2(new_n966), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT62), .B1(new_n996), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n966), .B1(new_n993), .B2(G286), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT51), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n995), .A4(new_n994), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT50), .B1(new_n988), .B2(new_n989), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .A3(new_n968), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n973), .B1(new_n969), .B2(new_n972), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n952), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n977), .A2(new_n973), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(new_n1012), .A3(new_n815), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n851), .A2(G1384), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n952), .B1(new_n1015), .B2(KEYINPUT45), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n694), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT55), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n697), .A2(G1976), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n969), .A2(new_n972), .A3(new_n968), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1027), .A2(new_n1028), .A3(G8), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1027), .B2(G8), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1024), .B(new_n1026), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G305), .B(G1981), .ZN(new_n1032));
  NOR2_X1   g607(.A1(KEYINPUT112), .A2(KEYINPUT49), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1032), .B(new_n1033), .Z(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1024), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT111), .B(new_n1024), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1018), .B1(G2090), .B2(new_n978), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1022), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(G8), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1023), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1017), .A2(G2078), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1047), .A2(new_n1048), .B1(new_n737), .B2(new_n978), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n985), .A2(new_n799), .A3(new_n986), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT53), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1046), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1003), .A2(new_n1007), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1035), .A2(new_n1025), .A3(new_n697), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(G1981), .B2(G305), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT113), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1042), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(new_n1045), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n993), .A2(G8), .A3(G168), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1046), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1066), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1043), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n1022), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n1045), .A3(new_n1042), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1064), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1057), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1027), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT110), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1027), .A2(new_n1028), .A3(G8), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(G1976), .B2(new_n697), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT52), .B1(new_n1078), .B2(KEYINPUT111), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1041), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1074), .B(new_n1045), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1044), .B1(new_n1019), .B2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(G171), .B(KEYINPUT54), .Z(new_n1084));
  NAND3_X1  g659(.A1(new_n799), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n480), .B(new_n1085), .C1(new_n1015), .C2(KEYINPUT45), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1086), .B2(new_n949), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1054), .A2(new_n1084), .B1(new_n1049), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1083), .B(new_n1088), .C1(new_n996), .C2(new_n1002), .ZN(new_n1089));
  XOR2_X1   g664(.A(G299), .B(KEYINPUT57), .Z(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1016), .B(new_n1092), .C1(new_n977), .C2(KEYINPUT45), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1091), .B1(new_n1097), .B2(KEYINPUT119), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1099), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT120), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n952), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(KEYINPUT114), .B1(new_n973), .B2(new_n977), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1956), .B1(new_n1103), .B2(new_n1012), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1099), .B1(new_n1104), .B2(new_n1094), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1091), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n978), .A2(new_n751), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1027), .A2(G2067), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT117), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(KEYINPUT117), .A3(new_n1110), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n614), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1112), .A2(KEYINPUT118), .A3(new_n614), .A4(new_n1113), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1101), .A2(new_n1108), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1097), .A2(new_n1090), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1093), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1124), .B2(new_n1091), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1119), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1113), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT60), .B(new_n606), .C1(new_n1128), .C2(new_n1111), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1027), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1017), .B2(G1996), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1132), .B(new_n560), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1132), .A2(new_n560), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n1134), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n1128), .B2(new_n1111), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1112), .A2(new_n1141), .A3(new_n1113), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1142), .A3(new_n614), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1097), .A2(KEYINPUT122), .A3(new_n1090), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1119), .B1(new_n1144), .B2(KEYINPUT61), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1127), .A2(new_n1139), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1089), .B1(new_n1120), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n963), .B1(new_n1073), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n953), .A2(new_n956), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT125), .ZN(new_n1152));
  INV_X1    g727(.A(new_n953), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n955), .B2(new_n854), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n714), .A2(new_n717), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n959), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n765), .A2(new_n954), .A3(new_n766), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G290), .A2(G1986), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n953), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n961), .A2(new_n953), .B1(KEYINPUT48), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(KEYINPUT48), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1161), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1157), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT126), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1148), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g745(.A(G319), .B1(new_n652), .B2(new_n653), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G227), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n689), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g748(.A(new_n1174), .B1(new_n944), .B2(new_n945), .ZN(new_n1175));
  AND3_X1   g749(.A1(new_n886), .A2(new_n1175), .A3(KEYINPUT127), .ZN(new_n1176));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n886), .B2(new_n1175), .ZN(new_n1177));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n1177), .ZN(G308));
  NAND2_X1  g752(.A1(new_n886), .A2(new_n1175), .ZN(G225));
endmodule


