//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G472), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT67), .A2(G131), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI211_X1 g008(.A(KEYINPUT66), .B(new_n193), .C1(new_n194), .C2(G137), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT66), .B1(new_n198), .B2(new_n193), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(G137), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n192), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n194), .A2(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(KEYINPUT11), .ZN(new_n207));
  AND4_X1   g021(.A1(new_n192), .A2(new_n203), .A3(new_n207), .A4(new_n195), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n191), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n192), .A3(new_n203), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n207), .A3(new_n195), .ZN(new_n211));
  INV_X1    g025(.A(new_n192), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT69), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT64), .A3(G143), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT0), .B(G128), .Z(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT0), .A3(G128), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n209), .A2(new_n214), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n216), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(G128), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n219), .A2(G143), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n218), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n198), .A2(new_n202), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n203), .A2(new_n207), .A3(new_n239), .A4(new_n195), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(KEYINPUT30), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT2), .B(G113), .Z(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n236), .A2(new_n247), .A3(new_n238), .A4(new_n240), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n223), .A2(new_n249), .A3(new_n225), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n223), .B2(new_n225), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n210), .A2(new_n213), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n246), .A2(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n242), .B(new_n245), .C1(KEYINPUT30), .C2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n245), .B(KEYINPUT70), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n227), .A2(new_n241), .A3(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n255), .A2(KEYINPUT31), .A3(new_n257), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n245), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n257), .B1(new_n269), .B2(new_n254), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n257), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n263), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n190), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n187), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n266), .A2(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n280), .C2(new_n190), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n255), .A2(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n275), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n284), .B(new_n285), .C1(new_n274), .C2(new_n275), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n227), .A2(new_n241), .ZN(new_n287));
  INV_X1    g101(.A(new_n256), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n272), .B1(new_n289), .B2(new_n257), .ZN(new_n290));
  INV_X1    g104(.A(new_n273), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n275), .A2(new_n285), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G140), .ZN(new_n299));
  XNOR2_X1  g113(.A(G125), .B(G140), .ZN(new_n300));
  MUX2_X1   g114(.A(new_n299), .B(new_n300), .S(KEYINPUT16), .Z(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(new_n219), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n232), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT24), .B(G110), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n303), .B1(KEYINPUT74), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n310), .B(new_n305), .C1(new_n311), .C2(new_n303), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G110), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n301), .A2(new_n219), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n300), .A2(new_n219), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(new_n307), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT75), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(new_n320), .C1(new_n312), .C2(G110), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n315), .B(new_n316), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n322), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT22), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(G137), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n314), .B(new_n329), .C1(new_n323), .C2(new_n324), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n189), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(G217), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(G217), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT73), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n331), .A2(new_n189), .A3(new_n334), .A4(new_n332), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n331), .A2(new_n332), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n340), .A2(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  XNOR2_X1  g164(.A(G104), .B(G107), .ZN(new_n351));
  INV_X1    g165(.A(G101), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT81), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n354), .B2(G107), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G104), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(G107), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n355), .A2(new_n358), .A3(new_n352), .A4(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n357), .A2(G104), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n354), .A2(G107), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n361), .B(G101), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n221), .A2(new_n230), .B1(new_n224), .B2(new_n233), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n232), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n235), .B1(new_n368), .B2(new_n224), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(new_n360), .A3(new_n364), .A4(new_n353), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n209), .A2(new_n371), .A3(new_n214), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT12), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n253), .A3(KEYINPUT12), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n374), .B2(new_n376), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n209), .A2(new_n214), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(G101), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n226), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n353), .A2(new_n360), .A3(new_n364), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT10), .A3(new_n236), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n379), .A2(new_n381), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G110), .B(G140), .Z(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT80), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n326), .A2(G227), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n377), .A2(new_n378), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n209), .A2(new_n214), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n387), .A3(new_n381), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(new_n390), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n350), .B(new_n189), .C1(new_n396), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n390), .A3(new_n394), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(new_n398), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n374), .B2(new_n376), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(G469), .C1(new_n404), .C2(new_n394), .ZN(new_n405));
  NAND2_X1  g219(.A1(G469), .A2(G902), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT9), .B(G234), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G221), .B1(new_n409), .B2(G902), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT79), .Z(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n232), .B2(G143), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n216), .A2(KEYINPUT93), .A3(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT13), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n232), .A2(G143), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n420), .A2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n194), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT94), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n427), .A2(KEYINPUT94), .ZN(new_n429));
  INV_X1    g243(.A(G116), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT92), .B1(new_n430), .B2(G122), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(G122), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(G107), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G107), .B1(new_n435), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n441));
  INV_X1    g255(.A(new_n427), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n194), .B1(new_n420), .B2(new_n423), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT95), .A3(new_n427), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n436), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT14), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n431), .B2(new_n434), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n449), .B2(new_n357), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n435), .A2(new_n448), .A3(G107), .A4(new_n436), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n440), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n409), .A2(new_n338), .A3(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n453), .A3(new_n455), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n189), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n461), .B(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n465));
  NOR2_X1   g279(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n466));
  OR3_X1    g280(.A1(new_n300), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n300), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n219), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n259), .A2(G214), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT89), .A3(G143), .ZN(new_n472));
  OR2_X1    g286(.A1(KEYINPUT89), .A2(G143), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT89), .A2(G143), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n473), .A2(G214), .A3(new_n259), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n239), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(G131), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n315), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n478), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT18), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n300), .B(new_n219), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n482), .A2(new_n484), .A3(new_n485), .A4(new_n477), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(G113), .B(G122), .Z(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT91), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n354), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n477), .A2(new_n493), .A3(new_n478), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n301), .A2(new_n219), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n481), .A2(KEYINPUT17), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n494), .A2(new_n315), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n490), .A3(new_n486), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G475), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n189), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n490), .B1(new_n497), .B2(new_n486), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n189), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G475), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n500), .A4(new_n189), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n464), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(G234), .A2(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G952), .A3(new_n326), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT97), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT21), .B(G898), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(G902), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n243), .A2(new_n244), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n523));
  OR3_X1    g337(.A1(new_n430), .A2(KEYINPUT5), .A3(G119), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(G113), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n388), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n245), .A2(new_n386), .A3(new_n384), .ZN(new_n527));
  XOR2_X1   g341(.A(G110), .B(G122), .Z(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n528), .B(KEYINPUT8), .Z(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n522), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(new_n365), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n365), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  INV_X1    g350(.A(G224), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT7), .B1(new_n537), .B2(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n366), .A2(G125), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n223), .A2(G125), .A3(new_n225), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n536), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  AND4_X1   g358(.A1(new_n530), .A2(new_n535), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT87), .B1(new_n543), .B2(new_n538), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n529), .B1(new_n526), .B2(new_n527), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n537), .A2(G953), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n543), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT85), .B(KEYINPUT6), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n548), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n548), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n550), .B(new_n552), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n547), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT88), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(new_n559), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT84), .Z(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n521), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n297), .A2(new_n349), .A3(new_n416), .A4(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G101), .ZN(G3));
  INV_X1    g384(.A(new_n277), .ZN(new_n571));
  OAI21_X1  g385(.A(G472), .B1(new_n280), .B2(G902), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n349), .A2(new_n416), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  INV_X1    g390(.A(new_n458), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n455), .B1(new_n440), .B2(new_n453), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n459), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n459), .B2(new_n576), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n457), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n458), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G478), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n459), .A2(new_n462), .A3(new_n189), .ZN(new_n589));
  NAND2_X1  g403(.A1(G478), .A2(G902), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n588), .A2(new_n509), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n565), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n559), .B1(new_n547), .B2(new_n557), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n594), .B2(new_n563), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n520), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n575), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT34), .B(G104), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  INV_X1    g414(.A(new_n509), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n464), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n575), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n325), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n344), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n342), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n607), .B1(new_n342), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n416), .A2(new_n568), .A3(new_n573), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT37), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G110), .ZN(G12));
  INV_X1    g430(.A(new_n563), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n565), .B1(new_n617), .B2(new_n593), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n413), .B2(new_n415), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n513), .B1(G900), .B2(new_n517), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n602), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n297), .A2(new_n619), .A3(new_n613), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G128), .ZN(G30));
  AND2_X1   g438(.A1(new_n289), .A2(new_n257), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n264), .B(G472), .C1(new_n263), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(G472), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT101), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n282), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n592), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n620), .B(KEYINPUT39), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n416), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n564), .B(KEYINPUT38), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n416), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n632), .A2(new_n635), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n613), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n464), .A2(new_n509), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n216), .ZN(G45));
  NOR2_X1   g458(.A1(new_n591), .A2(new_n621), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n297), .A2(new_n619), .A3(new_n613), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  NAND2_X1  g461(.A1(new_n374), .A2(new_n376), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT82), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n649), .A2(new_n390), .A3(new_n394), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n400), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n350), .B1(new_n653), .B2(new_n189), .ZN(new_n654));
  AOI211_X1 g468(.A(G469), .B(G902), .C1(new_n651), .C2(new_n652), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n410), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n297), .A2(new_n349), .A3(new_n597), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT41), .B(G113), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G15));
  NAND4_X1  g475(.A1(new_n297), .A2(new_n349), .A3(new_n603), .A4(new_n658), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G116), .ZN(G18));
  AOI21_X1  g477(.A(new_n188), .B1(new_n286), .B2(new_n294), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n279), .B2(new_n281), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n521), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n613), .A2(new_n410), .A3(new_n656), .A4(new_n595), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n665), .A2(new_n667), .A3(new_n670), .A4(new_n521), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n304), .ZN(G21));
  OAI21_X1  g487(.A(new_n275), .B1(new_n290), .B2(new_n291), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n190), .B1(new_n268), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n572), .A2(KEYINPUT103), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(G472), .C1(new_n280), .C2(G902), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n657), .A2(new_n519), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n641), .A2(new_n595), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n464), .A2(new_n509), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n618), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n679), .A2(new_n680), .A3(new_n346), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT105), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n433), .ZN(G24));
  NAND3_X1  g502(.A1(new_n668), .A2(new_n679), .A3(new_n645), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  AOI21_X1  g504(.A(new_n348), .B1(new_n282), .B2(new_n296), .ZN(new_n691));
  INV_X1    g505(.A(new_n591), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n620), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n405), .A2(KEYINPUT106), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n648), .A2(new_n390), .ZN(new_n696));
  INV_X1    g510(.A(new_n394), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n699), .A3(G469), .A4(new_n402), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n401), .A2(new_n695), .A3(new_n406), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT107), .A3(new_n410), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT107), .B1(new_n701), .B2(new_n410), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n564), .A2(new_n592), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n691), .A2(new_n694), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n187), .B1(new_n280), .B2(new_n190), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n296), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n645), .A3(new_n346), .A4(new_n705), .ZN(new_n712));
  INV_X1    g526(.A(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n702), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT42), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n239), .ZN(G33));
  INV_X1    g531(.A(new_n622), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n691), .A2(new_n707), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  OR2_X1    g536(.A1(new_n573), .A2(new_n640), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n573), .A2(new_n640), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n581), .A2(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n589), .B(new_n590), .C1(new_n728), .C2(new_n462), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  OR3_X1    g544(.A1(new_n729), .A2(new_n730), .A3(new_n509), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n729), .B2(new_n509), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n724), .A2(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n706), .B1(new_n736), .B2(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n698), .A2(new_n402), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n698), .A2(KEYINPUT45), .A3(new_n402), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(G469), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT46), .B1(new_n742), .B2(new_n406), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n655), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(KEYINPUT46), .A3(new_n406), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n410), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n633), .ZN(new_n749));
  INV_X1    g563(.A(new_n727), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n725), .A2(new_n726), .ZN(new_n751));
  INV_X1    g565(.A(new_n735), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n733), .A2(KEYINPUT109), .ZN(new_n753));
  OAI22_X1  g567(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n197), .ZN(G39));
  AND3_X1   g572(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n410), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT47), .B1(new_n746), .B2(new_n410), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n665), .B(new_n348), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n645), .A2(new_n705), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(G140), .Z(G42));
  NAND2_X1  g578(.A1(new_n701), .A2(new_n410), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n342), .A2(new_n610), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n682), .B2(new_n684), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n630), .A2(new_n620), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n623), .A2(new_n646), .A3(new_n769), .A4(new_n689), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n415), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n414), .B1(new_n407), .B2(new_n411), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n595), .B(new_n613), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n665), .A2(new_n718), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n665), .A2(new_n693), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(KEYINPUT52), .A3(new_n689), .A4(new_n769), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n519), .B(new_n567), .C1(new_n591), .C2(new_n602), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n349), .A3(new_n416), .A4(new_n573), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n569), .B(new_n785), .C1(new_n669), .C2(new_n671), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n721), .A2(new_n715), .A3(new_n708), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n659), .A2(new_n662), .A3(new_n614), .A4(new_n686), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n510), .A2(KEYINPUT111), .A3(new_n620), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT111), .B1(new_n510), .B2(new_n620), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n297), .A2(new_n416), .A3(new_n705), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n703), .A2(new_n704), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n679), .A3(new_n645), .A4(new_n705), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n640), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n772), .A2(KEYINPUT113), .A3(new_n780), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n783), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n772), .A2(new_n800), .A3(new_n780), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n569), .A2(new_n785), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n666), .A2(new_n668), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n670), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n666), .A2(KEYINPUT102), .A3(new_n668), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n787), .ZN(new_n808));
  INV_X1    g622(.A(new_n795), .ZN(new_n809));
  INV_X1    g623(.A(new_n788), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n800), .B1(new_n772), .B2(new_n780), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n802), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n799), .B1(new_n813), .B2(new_n797), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n657), .A2(new_n706), .A3(new_n513), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n631), .A2(new_n349), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n729), .A2(new_n601), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n679), .A2(new_n346), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n821), .A2(new_n514), .A3(new_n733), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n636), .A2(new_n657), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n592), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n592), .A3(new_n514), .A4(new_n733), .ZN(new_n827));
  INV_X1    g641(.A(new_n825), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT115), .B(new_n823), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n820), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n817), .A2(new_n733), .A3(KEYINPUT116), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT116), .B1(new_n817), .B2(new_n733), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n613), .B(new_n679), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n759), .A2(new_n760), .ZN(new_n834));
  INV_X1    g648(.A(new_n656), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(new_n411), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n705), .B(new_n822), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n830), .A2(KEYINPUT51), .A3(new_n833), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n822), .A2(new_n595), .A3(new_n658), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  INV_X1    g655(.A(G952), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n711), .A2(new_n346), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n831), .B2(new_n832), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT48), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT48), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n842), .B(G953), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n818), .A2(new_n692), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n839), .A2(new_n841), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n836), .B(KEYINPUT114), .Z(new_n851));
  OAI211_X1 g665(.A(new_n705), .B(new_n822), .C1(new_n834), .C2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n830), .A2(new_n833), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n783), .A2(new_n796), .A3(new_n798), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n781), .A2(KEYINPUT112), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n796), .A3(new_n797), .A4(new_n801), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n816), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n842), .A2(new_n326), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n816), .A2(new_n856), .A3(new_n861), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n411), .B1(new_n835), .B2(KEYINPUT49), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n868), .A2(new_n636), .A3(new_n509), .A4(new_n729), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n346), .A3(new_n566), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n631), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n872), .ZN(G75));
  NAND3_X1  g687(.A1(new_n859), .A2(new_n796), .A3(new_n801), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT53), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(G210), .A3(G902), .A4(new_n799), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n552), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT55), .Z(new_n881));
  AOI21_X1  g695(.A(KEYINPUT119), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  INV_X1    g697(.A(new_n881), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n883), .B(new_n884), .C1(new_n876), .C2(new_n877), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n326), .A2(G952), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n875), .A2(G902), .A3(new_n561), .A4(new_n799), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n886), .A2(new_n894), .ZN(G51));
  OR2_X1    g709(.A1(new_n406), .A2(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n406), .A2(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n875), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT54), .B1(new_n875), .B2(new_n799), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n896), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n653), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n875), .A2(G902), .A3(new_n799), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n742), .B(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n887), .B1(new_n902), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n498), .A3(new_n492), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .A4(new_n499), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(new_n888), .A3(new_n910), .ZN(G60));
  XOR2_X1   g725(.A(new_n590), .B(KEYINPUT59), .Z(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n728), .B(new_n913), .C1(new_n899), .C2(new_n900), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n816), .B2(new_n861), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n888), .C1(new_n728), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(G63));
  XOR2_X1   g731(.A(new_n337), .B(KEYINPUT60), .Z(new_n918));
  NAND4_X1  g732(.A1(new_n875), .A2(new_n609), .A3(new_n799), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n875), .A2(new_n799), .A3(new_n918), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n888), .B(new_n919), .C1(new_n921), .C2(new_n343), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G66));
  OAI21_X1  g738(.A(G953), .B1(new_n516), .B2(new_n537), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n786), .A2(new_n788), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n879), .B1(G898), .B2(new_n326), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  AOI21_X1  g743(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n779), .A2(new_n689), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n757), .A2(new_n932), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n843), .B(new_n749), .C1(new_n682), .C2(new_n684), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n934), .A2(new_n763), .A3(new_n787), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n326), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n242), .B1(KEYINPUT30), .B2(new_n254), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT122), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n469), .ZN(new_n939));
  NAND2_X1  g753(.A1(G900), .A2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n930), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n939), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n931), .B1(new_n642), .B2(new_n639), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n763), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n931), .B(new_n948), .C1(new_n642), .C2(new_n639), .ZN(new_n949));
  INV_X1    g763(.A(new_n602), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n691), .B1(new_n692), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n951), .A2(new_n634), .A3(new_n706), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n737), .B2(new_n756), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n947), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n944), .B1(new_n954), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n943), .B(new_n956), .Z(G72));
  NAND4_X1  g771(.A1(new_n947), .A2(new_n926), .A3(new_n953), .A4(new_n949), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n627), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n275), .B1(new_n961), .B2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n958), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n283), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n284), .A2(new_n264), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n858), .A2(new_n860), .A3(new_n960), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n888), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n933), .A2(new_n926), .A3(new_n935), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n263), .B(new_n283), .C1(new_n971), .C2(new_n960), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(G57));
endmodule


