//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT79), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT80), .A4(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G101), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(KEYINPUT81), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n213), .A2(new_n219), .A3(G101), .A4(new_n214), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n206), .A2(new_n209), .A3(new_n221), .A4(new_n210), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AND4_X1   g038(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n215), .B2(KEYINPUT81), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n217), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n204), .B(new_n216), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G128), .A3(new_n202), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n195), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(new_n202), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n210), .A2(KEYINPUT83), .ZN(new_n237));
  INV_X1    g051(.A(new_n210), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT83), .B1(new_n205), .B2(G107), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(G101), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n222), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n235), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n240), .A2(new_n222), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT84), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n229), .A2(KEYINPUT84), .A3(G128), .A4(new_n202), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n231), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT85), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n202), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n243), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n242), .B1(new_n236), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n228), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT87), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT64), .B1(new_n260), .B2(G134), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n258), .B2(G137), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT11), .ZN(new_n266));
  OAI21_X1  g080(.A(G131), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n260), .A2(G134), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n265), .B2(KEYINPUT11), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n261), .A2(new_n262), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT65), .B(G131), .C1(new_n263), .C2(new_n266), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n228), .A2(new_n255), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n257), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n276), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n228), .A2(new_n255), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n193), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n193), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT86), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n235), .A2(new_n241), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n254), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  AND4_X1   g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n276), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n284), .A2(new_n287), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT86), .A2(KEYINPUT12), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n289), .B(new_n290), .C1(new_n286), .C2(new_n276), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n283), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n187), .B(new_n188), .C1(new_n282), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(G469), .A2(G902), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n291), .A2(new_n288), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  INV_X1    g110(.A(new_n193), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n279), .ZN(new_n299));
  OAI211_X1 g113(.A(G469), .B(new_n298), .C1(new_n299), .C2(new_n283), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT78), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G110), .B(G122), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT2), .B(G113), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n216), .C1(new_n225), .C2(new_n227), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n311), .A2(new_n312), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT5), .ZN(new_n317));
  OAI21_X1  g131(.A(G113), .B1(new_n308), .B2(KEYINPUT5), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n243), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n306), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT6), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT6), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n321), .A3(new_n306), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n315), .A2(KEYINPUT88), .A3(new_n321), .A4(new_n306), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n323), .B1(new_n329), .B2(new_n322), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n235), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n331), .B2(new_n204), .ZN(new_n333));
  INV_X1    g147(.A(G224), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT7), .B1(new_n334), .B2(G953), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n333), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n306), .B(KEYINPUT8), .Z(new_n340));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n318), .B1(new_n317), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n341), .B2(new_n317), .ZN(new_n343));
  INV_X1    g157(.A(new_n316), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n241), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n340), .B(new_n345), .C1(new_n241), .C2(new_n320), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n346), .A2(KEYINPUT90), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(KEYINPUT90), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n339), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n327), .A2(new_n328), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G210), .B1(G237), .B2(G902), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n353), .B(KEYINPUT91), .Z(new_n354));
  XOR2_X1   g168(.A(new_n354), .B(KEYINPUT92), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n354), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n337), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G128), .B(G143), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n258), .ZN(new_n361));
  XNOR2_X1  g175(.A(G116), .B(G122), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n208), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n309), .A2(KEYINPUT14), .A3(G122), .ZN(new_n364));
  XOR2_X1   g178(.A(G116), .B(G122), .Z(new_n365));
  OAI211_X1 g179(.A(G107), .B(new_n364), .C1(new_n365), .C2(KEYINPUT14), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n363), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n258), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n231), .A2(KEYINPUT13), .A3(G143), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n258), .B(new_n372), .C1(KEYINPUT13), .C2(new_n360), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n367), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n303), .A2(new_n375), .A3(G953), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n374), .B(new_n376), .Z(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(new_n188), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT15), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G478), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(KEYINPUT97), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(KEYINPUT97), .A3(new_n188), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n379), .A3(G478), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n381), .A2(KEYINPUT98), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT98), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n205), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  AOI21_X1  g205(.A(G140), .B1(new_n391), .B2(KEYINPUT75), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT75), .B1(new_n331), .B2(KEYINPUT74), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(G140), .B2(new_n396), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n397), .A2(KEYINPUT94), .A3(new_n194), .ZN(new_n398));
  INV_X1    g212(.A(G237), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT68), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT68), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G237), .ZN(new_n402));
  AOI21_X1  g216(.A(G953), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT93), .B(G143), .Z(new_n404));
  AND3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(G214), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n196), .A2(KEYINPUT93), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n403), .B2(G214), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT18), .B(G131), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n403), .A2(new_n404), .A3(G214), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n194), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT94), .B(new_n414), .C1(new_n397), .C2(new_n194), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n398), .A2(new_n408), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G140), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT16), .B1(new_n417), .B2(G125), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT16), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n397), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G146), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n194), .B(new_n419), .C1(new_n397), .C2(new_n420), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(new_n271), .A3(new_n411), .ZN(new_n424));
  OAI21_X1  g238(.A(G131), .B1(new_n405), .B2(new_n407), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n422), .B(new_n423), .C1(new_n426), .C2(KEYINPUT17), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT17), .B(G131), .C1(new_n405), .C2(new_n407), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n389), .B(new_n416), .C1(new_n427), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n422), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n413), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n397), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G146), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n416), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n389), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT96), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n440), .A2(new_n445), .A3(new_n441), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT20), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n427), .A2(new_n430), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n389), .B1(new_n450), .B2(new_n416), .ZN(new_n451));
  INV_X1    g265(.A(new_n431), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n188), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G475), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G952), .ZN(new_n458));
  AOI211_X1 g272(.A(G953), .B(new_n458), .C1(G234), .C2(G237), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT99), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n188), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR4_X1   g278(.A1(new_n387), .A2(new_n455), .A3(new_n457), .A4(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(G119), .B(G128), .Z(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT24), .B(G110), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT73), .B1(new_n307), .B2(G128), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n473), .A2(KEYINPUT23), .B1(new_n307), .B2(G128), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(KEYINPUT23), .B2(new_n473), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n475), .B2(G110), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n422), .A2(new_n414), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n475), .B2(G110), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n423), .B2(new_n422), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n469), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n422), .A2(new_n423), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n479), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n422), .A2(new_n414), .A3(new_n476), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n468), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n486), .A3(new_n188), .ZN(new_n487));
  NOR2_X1   g301(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n482), .A2(new_n486), .A3(new_n188), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n375), .B1(G234), .B2(new_n188), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n482), .A2(new_n486), .ZN(new_n495));
  INV_X1    g309(.A(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n188), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT77), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n274), .A2(new_n275), .A3(new_n204), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n258), .A2(G137), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n506), .B2(new_n269), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n234), .A2(new_n273), .A3(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n505), .A2(new_n501), .A3(new_n502), .A4(new_n508), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n314), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n403), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n313), .A3(new_n508), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n505), .A2(new_n508), .ZN(new_n523));
  INV_X1    g337(.A(new_n503), .ZN(new_n524));
  INV_X1    g338(.A(new_n504), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n510), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n522), .B1(new_n527), .B2(new_n314), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT31), .A3(new_n517), .ZN(new_n529));
  INV_X1    g343(.A(new_n517), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n522), .A2(KEYINPUT28), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n314), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(new_n518), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n531), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n521), .A2(new_n529), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(G472), .A2(G902), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT32), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n530), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT31), .B1(new_n528), .B2(new_n517), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n313), .B1(new_n526), .B2(new_n510), .ZN(new_n544));
  NOR4_X1   g358(.A1(new_n544), .A2(new_n530), .A3(new_n520), .A4(new_n522), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n539), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n537), .A2(new_n530), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n530), .B1(new_n544), .B2(new_n522), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n550), .A2(KEYINPUT29), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n532), .A2(new_n554), .A3(new_n518), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n314), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(KEYINPUT28), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n531), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n517), .A2(KEYINPUT29), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n188), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G472), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n500), .B1(new_n549), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n305), .A2(new_n359), .A3(new_n465), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  OAI21_X1  g378(.A(G472), .B1(new_n538), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n546), .A2(new_n539), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n500), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n305), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n570));
  INV_X1    g384(.A(new_n464), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n337), .A2(new_n351), .A3(new_n357), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n357), .B1(new_n337), .B2(new_n351), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n456), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G478), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n378), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n188), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n377), .B(KEYINPUT33), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n576), .B(new_n578), .C1(new_n579), .C2(new_n575), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n455), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n570), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n352), .A2(new_n354), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n457), .B1(new_n584), .B2(new_n358), .ZN(new_n585));
  INV_X1    g399(.A(new_n582), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(KEYINPUT100), .A3(new_n571), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n569), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT102), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NAND2_X1  g406(.A1(new_n448), .A2(new_n443), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n454), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n569), .A2(new_n574), .A3(new_n386), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT35), .B(G107), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G9));
  NAND2_X1  g411(.A1(new_n484), .A2(new_n485), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT103), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n598), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n498), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n494), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT104), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n492), .A2(new_n493), .B1(new_n498), .B2(new_n601), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n567), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n305), .A2(new_n359), .A3(new_n465), .A4(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT37), .B(G110), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  NOR3_X1   g426(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n547), .B1(new_n546), .B2(new_n539), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n561), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n615), .A2(new_n304), .A3(new_n301), .ZN(new_n616));
  INV_X1    g430(.A(new_n608), .ZN(new_n617));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n459), .B1(new_n463), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n386), .A2(new_n594), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n585), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G128), .ZN(G30));
  XOR2_X1   g436(.A(new_n619), .B(KEYINPUT39), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n305), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n359), .A2(KEYINPUT38), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n356), .A2(new_n628), .A3(new_n358), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n555), .A2(new_n530), .A3(new_n556), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(KEYINPUT105), .ZN(new_n632));
  INV_X1    g446(.A(new_n519), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(KEYINPUT105), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n549), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n549), .A2(KEYINPUT106), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n449), .A2(new_n454), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n386), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n456), .A2(new_n641), .A3(new_n605), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n626), .A2(new_n630), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G143), .ZN(G45));
  AOI211_X1 g460(.A(new_n619), .B(new_n580), .C1(new_n449), .C2(new_n454), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n616), .A2(new_n585), .A3(new_n617), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  NAND2_X1  g463(.A1(new_n279), .A2(new_n281), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n292), .B1(new_n650), .B2(new_n297), .ZN(new_n651));
  OAI21_X1  g465(.A(G469), .B1(new_n651), .B2(G902), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n304), .A3(new_n293), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n562), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n583), .B2(new_n587), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT41), .B(G113), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G15));
  OAI21_X1  g472(.A(new_n456), .B1(new_n572), .B2(new_n573), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n660), .A2(new_n615), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n494), .A2(new_n499), .A3(new_n571), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n386), .A2(new_n594), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  NOR4_X1   g479(.A1(new_n608), .A2(new_n387), .A3(new_n455), .A4(new_n464), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  INV_X1    g482(.A(G472), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n546), .B2(new_n188), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n521), .A2(new_n529), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n558), .A2(new_n530), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n540), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OR3_X1    g487(.A1(new_n670), .A2(new_n662), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n653), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n585), .A3(KEYINPUT107), .A4(new_n643), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n456), .B(new_n643), .C1(new_n572), .C2(new_n573), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n670), .A2(new_n662), .A3(new_n673), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n304), .A3(new_n293), .A4(new_n652), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G122), .ZN(G24));
  INV_X1    g497(.A(new_n673), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n565), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n605), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n585), .A2(new_n654), .A3(new_n647), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G125), .ZN(G27));
  INV_X1    g502(.A(new_n355), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n337), .B2(new_n351), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n572), .A2(new_n690), .A3(new_n457), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n294), .B(KEYINPUT108), .Z(new_n692));
  NAND3_X1  g506(.A1(new_n293), .A2(new_n300), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n304), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n691), .A2(new_n695), .A3(new_n562), .A4(new_n647), .ZN(new_n696));
  NOR2_X1   g510(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n356), .A2(new_n358), .A3(new_n456), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n694), .ZN(new_n700));
  INV_X1    g514(.A(new_n697), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n562), .A3(new_n647), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n562), .A3(new_n620), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G134), .ZN(G36));
  NAND2_X1  g520(.A1(new_n567), .A2(new_n603), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT112), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n455), .A2(KEYINPUT43), .A3(new_n580), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n642), .A2(KEYINPUT111), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n455), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n581), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n713), .B2(KEYINPUT43), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT44), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n699), .ZN(new_n716));
  OAI211_X1 g530(.A(KEYINPUT45), .B(new_n298), .C1(new_n299), .C2(new_n283), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n280), .B1(new_n256), .B2(KEYINPUT87), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n283), .B1(new_n719), .B2(new_n278), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n193), .B1(new_n295), .B2(new_n281), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n722), .A3(G469), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n692), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n293), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n304), .B(new_n623), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n708), .A2(KEYINPUT44), .A3(new_n714), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n716), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  OAI21_X1  g548(.A(new_n304), .B1(new_n727), .B2(new_n728), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(KEYINPUT47), .B(new_n304), .C1(new_n727), .C2(new_n728), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n647), .A2(new_n500), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n699), .A2(new_n615), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  NAND2_X1  g557(.A1(new_n458), .A2(new_n189), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n745));
  INV_X1    g559(.A(new_n459), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n685), .A2(new_n500), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n714), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n653), .A2(new_n456), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n627), .A2(new_n629), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT116), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n627), .A2(new_n752), .A3(new_n629), .A4(new_n749), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n641), .A2(new_n500), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n699), .A2(new_n746), .A3(new_n653), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n455), .A2(new_n581), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n686), .A3(new_n714), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n754), .B2(new_n755), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT117), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n652), .A2(new_n293), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n304), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n737), .A2(new_n738), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n748), .A2(new_n699), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n757), .A2(new_n764), .A3(KEYINPUT117), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n745), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n758), .A2(new_n586), .A3(new_n759), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n458), .A2(G953), .ZN(new_n777));
  INV_X1    g591(.A(new_n660), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n748), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT119), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT119), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n759), .A2(new_n562), .A3(new_n714), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT48), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n751), .A2(new_n753), .ZN(new_n785));
  INV_X1    g599(.A(new_n748), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n745), .B1(new_n770), .B2(new_n771), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n756), .A4(new_n763), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT118), .ZN(new_n791));
  INV_X1    g605(.A(new_n764), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n756), .A4(new_n789), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n784), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n775), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n621), .A2(new_n648), .A3(new_n687), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n603), .A2(new_n619), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n639), .B2(new_n640), .ZN(new_n800));
  INV_X1    g614(.A(new_n678), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n800), .A2(new_n801), .A3(new_n695), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n797), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n617), .B(new_n456), .C1(new_n572), .C2(new_n573), .ZN(new_n804));
  INV_X1    g618(.A(new_n620), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n615), .A2(new_n301), .A3(new_n304), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n647), .A2(new_n565), .A3(new_n603), .A4(new_n684), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n659), .A2(new_n808), .A3(new_n653), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n800), .A2(new_n801), .A3(new_n695), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(KEYINPUT52), .A3(new_n648), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n803), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n660), .B(new_n615), .C1(new_n663), .C2(new_n666), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n682), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n571), .A2(new_n456), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n381), .A2(new_n383), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n449), .A2(new_n454), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n582), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n305), .A2(new_n359), .A3(new_n568), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n563), .A2(new_n610), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n815), .A2(new_n656), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n699), .A2(new_n808), .A3(new_n694), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n594), .A2(new_n817), .A3(new_n619), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n699), .A2(new_n608), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n616), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n703), .A2(new_n705), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n813), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n583), .A2(new_n587), .ZN(new_n831));
  INV_X1    g645(.A(new_n655), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n821), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n682), .A4(new_n814), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n703), .A2(new_n705), .A3(new_n826), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n837), .B2(new_n813), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n828), .A2(new_n829), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT114), .B1(new_n815), .B2(new_n656), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n833), .A2(new_n845), .A3(new_n682), .A4(new_n814), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n813), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n840), .A2(new_n841), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n744), .B1(new_n796), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n713), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n766), .A2(KEYINPUT49), .ZN(new_n852));
  INV_X1    g666(.A(new_n304), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n500), .A2(new_n853), .A3(new_n457), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n766), .A2(KEYINPUT49), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n630), .A2(new_n855), .A3(new_n641), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT113), .Z(new_n858));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n858), .ZN(G75));
  XNOR2_X1  g673(.A(new_n330), .B(new_n336), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT55), .Z(new_n861));
  AOI21_X1  g675(.A(new_n188), .B1(new_n840), .B2(new_n847), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n354), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n864), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n862), .B2(new_n355), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n189), .A2(G952), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT120), .Z(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n865), .A2(new_n867), .A3(new_n870), .ZN(G51));
  XOR2_X1   g685(.A(new_n692), .B(KEYINPUT57), .Z(new_n872));
  AND3_X1   g686(.A1(new_n840), .A2(new_n841), .A3(new_n847), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n841), .B1(new_n840), .B2(new_n847), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n651), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n840), .A2(new_n847), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(G902), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(new_n723), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n868), .B1(new_n877), .B2(new_n880), .ZN(G54));
  NAND2_X1  g695(.A1(KEYINPUT58), .A2(G475), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n431), .B(new_n439), .C1(new_n879), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n868), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .A4(new_n440), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G60));
  XNOR2_X1  g700(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n578), .B(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n579), .B(new_n888), .C1(new_n873), .C2(new_n874), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n869), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n579), .B1(new_n849), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(G63));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n893));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT60), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n840), .B2(new_n847), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n601), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n869), .B1(new_n896), .B2(new_n495), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n495), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n840), .A2(new_n847), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n895), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT61), .A3(new_n869), .A4(new_n897), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n904), .ZN(G66));
  AOI21_X1  g719(.A(new_n189), .B1(new_n461), .B2(G224), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT122), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n822), .B2(G953), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT123), .Z(new_n909));
  OAI221_X1 g723(.A(new_n323), .B1(G898), .B2(new_n189), .C1(new_n329), .C2(new_n322), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(G69));
  NAND2_X1  g725(.A1(new_n618), .A2(G953), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n730), .A2(new_n562), .A3(new_n801), .A4(new_n731), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n703), .A3(new_n705), .A4(new_n742), .ZN(new_n914));
  INV_X1    g728(.A(new_n798), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n733), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n733), .A2(KEYINPUT125), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n527), .B(new_n435), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n189), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n912), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n645), .A2(new_n915), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n645), .A2(KEYINPUT62), .A3(new_n915), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n562), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n582), .A2(new_n818), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n624), .A2(new_n930), .A3(new_n699), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n733), .A2(new_n934), .A3(new_n742), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n922), .B1(new_n936), .B2(new_n189), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n924), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n924), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G72));
  NAND2_X1  g757(.A1(new_n528), .A2(new_n530), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n920), .A2(new_n822), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n929), .A2(new_n935), .A3(new_n822), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n530), .B(new_n528), .C1(new_n949), .C2(new_n947), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n830), .A2(new_n838), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n552), .B2(new_n633), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n884), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n948), .A2(new_n950), .A3(new_n953), .ZN(G57));
endmodule


