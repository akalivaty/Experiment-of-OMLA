

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753;

  AND2_X1 U369 ( .A1(n350), .A2(n349), .ZN(n432) );
  INV_X1 U370 ( .A(n721), .ZN(n349) );
  AND2_X1 U371 ( .A1(n429), .A2(n428), .ZN(n619) );
  NOR2_X1 U372 ( .A1(n617), .A2(n750), .ZN(n618) );
  XNOR2_X1 U373 ( .A(n568), .B(n427), .ZN(n371) );
  AND2_X1 U374 ( .A1(n404), .A2(n358), .ZN(n566) );
  XNOR2_X1 U375 ( .A(n376), .B(n375), .ZN(n404) );
  NOR2_X1 U376 ( .A1(n352), .A2(n596), .ZN(n604) );
  BUF_X1 U377 ( .A(n352), .Z(n347) );
  INV_X1 U378 ( .A(n592), .ZN(n352) );
  XNOR2_X1 U379 ( .A(n601), .B(n361), .ZN(n674) );
  XNOR2_X1 U380 ( .A(n523), .B(n424), .ZN(n558) );
  XNOR2_X1 U381 ( .A(n543), .B(n486), .ZN(n402) );
  INV_X1 U382 ( .A(KEYINPUT3), .ZN(n422) );
  INV_X1 U383 ( .A(G125), .ZN(n417) );
  INV_X2 U384 ( .A(G128), .ZN(n485) );
  NAND2_X1 U385 ( .A1(n348), .A2(n601), .ZN(n611) );
  XNOR2_X1 U386 ( .A(n599), .B(n598), .ZN(n348) );
  XNOR2_X1 U387 ( .A(n641), .B(n351), .ZN(n350) );
  INV_X1 U388 ( .A(n640), .ZN(n351) );
  XNOR2_X2 U389 ( .A(n422), .B(G119), .ZN(n416) );
  AND2_X1 U390 ( .A1(n476), .A2(n644), .ZN(n415) );
  AND2_X2 U391 ( .A1(n410), .A2(n411), .ZN(n379) );
  OR2_X2 U392 ( .A1(n365), .A2(n457), .ZN(n633) );
  XNOR2_X2 U393 ( .A(n498), .B(n497), .ZN(n601) );
  XNOR2_X2 U394 ( .A(n503), .B(n502), .ZN(n592) );
  NAND2_X1 U395 ( .A1(n413), .A2(n446), .ZN(n445) );
  OR2_X1 U396 ( .A1(n748), .A2(n397), .ZN(n393) );
  XNOR2_X1 U397 ( .A(n456), .B(KEYINPUT40), .ZN(n748) );
  AND2_X1 U398 ( .A1(n620), .A2(n660), .ZN(n456) );
  OR2_X1 U399 ( .A1(n573), .A2(n360), .ZN(n448) );
  XNOR2_X1 U400 ( .A(n389), .B(KEYINPUT75), .ZN(n613) );
  XNOR2_X1 U401 ( .A(n518), .B(KEYINPUT33), .ZN(n682) );
  AND2_X1 U402 ( .A1(n576), .A2(n577), .ZN(n660) );
  XOR2_X1 U403 ( .A(G137), .B(G140), .Z(n490) );
  OR2_X1 U404 ( .A1(n365), .A2(n459), .ZN(n716) );
  OR2_X1 U405 ( .A1(n365), .A2(n460), .ZN(n709) );
  OR2_X1 U406 ( .A1(n365), .A2(n458), .ZN(n641) );
  NAND2_X1 U407 ( .A1(n369), .A2(n366), .ZN(n582) );
  XNOR2_X1 U408 ( .A(n489), .B(n488), .ZN(n732) );
  AND2_X1 U409 ( .A1(n463), .A2(n387), .ZN(n386) );
  NAND2_X1 U410 ( .A1(n393), .A2(n392), .ZN(n396) );
  NOR2_X1 U411 ( .A1(n711), .A2(G902), .ZN(n498) );
  OR2_X1 U412 ( .A1(n639), .A2(G902), .ZN(n399) );
  INV_X1 U413 ( .A(KEYINPUT10), .ZN(n424) );
  XOR2_X1 U414 ( .A(G902), .B(KEYINPUT15), .Z(n526) );
  NAND2_X1 U415 ( .A1(n386), .A2(n672), .ZN(n381) );
  XOR2_X1 U416 ( .A(KEYINPUT97), .B(n580), .Z(n689) );
  NAND2_X1 U417 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U418 ( .A1(n412), .A2(KEYINPUT44), .ZN(n408) );
  NAND2_X1 U419 ( .A1(n584), .A2(n583), .ZN(n446) );
  XNOR2_X1 U420 ( .A(n581), .B(n378), .ZN(n584) );
  INV_X1 U421 ( .A(KEYINPUT65), .ZN(n378) );
  AND2_X1 U422 ( .A1(n396), .A2(n394), .ZN(n428) );
  NAND2_X1 U423 ( .A1(n674), .A2(n673), .ZN(n570) );
  NAND2_X1 U424 ( .A1(n352), .A2(n461), .ZN(n391) );
  INV_X1 U425 ( .A(n595), .ZN(n461) );
  XNOR2_X1 U426 ( .A(n732), .B(n400), .ZN(n639) );
  XNOR2_X1 U427 ( .A(n515), .B(n462), .ZN(n400) );
  XNOR2_X1 U428 ( .A(n507), .B(n508), .ZN(n462) );
  XNOR2_X1 U429 ( .A(G128), .B(KEYINPUT77), .ZN(n477) );
  XNOR2_X1 U430 ( .A(n480), .B(n421), .ZN(n420) );
  INV_X1 U431 ( .A(KEYINPUT89), .ZN(n421) );
  XNOR2_X1 U432 ( .A(G119), .B(G110), .ZN(n480) );
  XNOR2_X1 U433 ( .A(n558), .B(n423), .ZN(n736) );
  INV_X1 U434 ( .A(n490), .ZN(n423) );
  XNOR2_X1 U435 ( .A(n545), .B(n356), .ZN(n418) );
  XNOR2_X1 U436 ( .A(G122), .B(G134), .ZN(n540) );
  XNOR2_X1 U437 ( .A(n732), .B(n452), .ZN(n711) );
  XNOR2_X1 U438 ( .A(n453), .B(n495), .ZN(n452) );
  XNOR2_X1 U439 ( .A(n493), .B(n374), .ZN(n453) );
  NOR2_X1 U440 ( .A1(n688), .A2(n687), .ZN(n594) );
  AND2_X1 U441 ( .A1(n597), .A2(n604), .ZN(n599) );
  XNOR2_X1 U442 ( .A(n443), .B(n440), .ZN(n714) );
  XNOR2_X1 U443 ( .A(n555), .B(n441), .ZN(n440) );
  XNOR2_X1 U444 ( .A(n556), .B(n442), .ZN(n441) );
  NAND2_X1 U445 ( .A1(n526), .A2(G475), .ZN(n459) );
  NOR2_X1 U446 ( .A1(G952), .A2(n722), .ZN(n721) );
  NAND2_X1 U447 ( .A1(n689), .A2(KEYINPUT98), .ZN(n383) );
  AND2_X1 U448 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U449 ( .A1(n751), .A2(KEYINPUT82), .ZN(n368) );
  NAND2_X1 U450 ( .A1(n435), .A2(KEYINPUT47), .ZN(n434) );
  XOR2_X1 U451 ( .A(G137), .B(KEYINPUT5), .Z(n512) );
  XNOR2_X1 U452 ( .A(G116), .B(KEYINPUT92), .ZN(n509) );
  XOR2_X1 U453 ( .A(KEYINPUT93), .B(KEYINPUT74), .Z(n510) );
  INV_X1 U454 ( .A(G146), .ZN(n506) );
  XNOR2_X1 U455 ( .A(G101), .B(G113), .ZN(n508) );
  XOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n541) );
  XNOR2_X1 U457 ( .A(G131), .B(KEYINPUT67), .ZN(n487) );
  NOR2_X1 U458 ( .A1(G953), .A2(G237), .ZN(n552) );
  XNOR2_X1 U459 ( .A(n496), .B(n492), .ZN(n374) );
  XNOR2_X1 U460 ( .A(n491), .B(G146), .ZN(n492) );
  INV_X1 U461 ( .A(G107), .ZN(n491) );
  OR2_X1 U462 ( .A1(G902), .A2(G237), .ZN(n529) );
  XNOR2_X1 U463 ( .A(n431), .B(n373), .ZN(n684) );
  XNOR2_X1 U464 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n373) );
  AND2_X1 U465 ( .A1(n573), .A2(n360), .ZN(n450) );
  AND2_X1 U466 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U467 ( .A(G110), .B(G101), .Z(n520) );
  XNOR2_X1 U468 ( .A(n519), .B(G113), .ZN(n551) );
  XNOR2_X1 U469 ( .A(G104), .B(G122), .ZN(n519) );
  XNOR2_X1 U470 ( .A(G140), .B(G143), .ZN(n556) );
  INV_X1 U471 ( .A(KEYINPUT94), .ZN(n442) );
  INV_X1 U472 ( .A(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U473 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U474 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n522) );
  INV_X1 U475 ( .A(KEYINPUT84), .ZN(n521) );
  INV_X1 U476 ( .A(KEYINPUT45), .ZN(n444) );
  XNOR2_X1 U477 ( .A(n622), .B(n426), .ZN(n425) );
  INV_X1 U478 ( .A(KEYINPUT105), .ZN(n426) );
  INV_X1 U479 ( .A(KEYINPUT22), .ZN(n375) );
  NOR2_X1 U480 ( .A1(n672), .A2(n570), .ZN(n679) );
  BUF_X1 U481 ( .A(n625), .Z(n431) );
  NAND2_X1 U482 ( .A1(n390), .A2(n377), .ZN(n389) );
  NOR2_X1 U483 ( .A1(n391), .A2(n591), .ZN(n390) );
  INV_X1 U484 ( .A(KEYINPUT19), .ZN(n530) );
  INV_X1 U485 ( .A(KEYINPUT100), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n560), .B(n559), .ZN(n577) );
  OR2_X1 U487 ( .A1(n575), .A2(n597), .ZN(n464) );
  XNOR2_X1 U488 ( .A(n597), .B(n516), .ZN(n603) );
  XNOR2_X1 U489 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n516) );
  NAND2_X1 U490 ( .A1(n404), .A2(n403), .ZN(n568) );
  NAND2_X1 U491 ( .A1(n526), .A2(G472), .ZN(n458) );
  XNOR2_X1 U492 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U493 ( .A(n469), .B(n468), .ZN(n401) );
  XNOR2_X1 U494 ( .A(n542), .B(n520), .ZN(n468) );
  XNOR2_X1 U495 ( .A(n470), .B(n551), .ZN(n469) );
  XNOR2_X1 U496 ( .A(n416), .B(KEYINPUT16), .ZN(n470) );
  NAND2_X1 U497 ( .A1(n526), .A2(G217), .ZN(n457) );
  XNOR2_X1 U498 ( .A(n479), .B(n420), .ZN(n481) );
  XNOR2_X1 U499 ( .A(n544), .B(n418), .ZN(n548) );
  XNOR2_X1 U500 ( .A(n471), .B(n401), .ZN(n707) );
  XNOR2_X1 U501 ( .A(n473), .B(n472), .ZN(n471) );
  XNOR2_X1 U502 ( .A(n525), .B(n521), .ZN(n472) );
  XNOR2_X1 U503 ( .A(n402), .B(n524), .ZN(n473) );
  NAND2_X1 U504 ( .A1(n526), .A2(G210), .ZN(n460) );
  XNOR2_X1 U505 ( .A(n602), .B(KEYINPUT42), .ZN(n752) );
  NAND2_X1 U506 ( .A1(n371), .A2(n355), .ZN(n567) );
  XNOR2_X1 U507 ( .A(n714), .B(n474), .ZN(n715) );
  XNOR2_X1 U508 ( .A(n467), .B(n466), .ZN(n465) );
  XNOR2_X1 U509 ( .A(n711), .B(n364), .ZN(n466) );
  AND2_X1 U510 ( .A1(n704), .A2(n419), .ZN(n705) );
  AND2_X1 U511 ( .A1(n703), .A2(n722), .ZN(n419) );
  INV_X1 U512 ( .A(n674), .ZN(n403) );
  AND2_X1 U513 ( .A1(n448), .A2(n615), .ZN(n353) );
  NOR2_X1 U514 ( .A1(n365), .A2(n632), .ZN(n354) );
  NOR2_X1 U515 ( .A1(n347), .A2(n597), .ZN(n355) );
  XNOR2_X1 U516 ( .A(n593), .B(KEYINPUT39), .ZN(n620) );
  XNOR2_X1 U517 ( .A(KEYINPUT95), .B(KEYINPUT7), .ZN(n356) );
  AND2_X1 U518 ( .A1(n382), .A2(n385), .ZN(n357) );
  INV_X1 U519 ( .A(n689), .ZN(n463) );
  AND2_X1 U520 ( .A1(n475), .A2(n674), .ZN(n358) );
  AND2_X1 U521 ( .A1(n355), .A2(KEYINPUT82), .ZN(n359) );
  XNOR2_X1 U522 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n360) );
  XNOR2_X1 U523 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n361) );
  XOR2_X1 U524 ( .A(KEYINPUT102), .B(KEYINPUT30), .Z(n362) );
  AND2_X1 U525 ( .A1(KEYINPUT44), .A2(n414), .ZN(n363) );
  INV_X1 U526 ( .A(KEYINPUT80), .ZN(n414) );
  INV_X1 U527 ( .A(KEYINPUT98), .ZN(n387) );
  XOR2_X1 U528 ( .A(n713), .B(n712), .Z(n364) );
  INV_X1 U529 ( .A(G953), .ZN(n722) );
  XNOR2_X1 U530 ( .A(n365), .B(KEYINPUT78), .ZN(n704) );
  XNOR2_X2 U531 ( .A(n631), .B(KEYINPUT2), .ZN(n365) );
  NAND2_X1 U532 ( .A1(n371), .A2(n359), .ZN(n367) );
  NAND2_X1 U533 ( .A1(n370), .A2(n567), .ZN(n369) );
  NOR2_X1 U534 ( .A1(n751), .A2(KEYINPUT82), .ZN(n370) );
  XNOR2_X2 U535 ( .A(n566), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U536 ( .A1(n372), .A2(n565), .ZN(n376) );
  NAND2_X1 U537 ( .A1(n679), .A2(n372), .ZN(n571) );
  XNOR2_X1 U538 ( .A(n372), .B(n539), .ZN(n573) );
  XNOR2_X2 U539 ( .A(n538), .B(KEYINPUT0), .ZN(n372) );
  OR2_X2 U540 ( .A1(n582), .A2(n749), .ZN(n412) );
  XNOR2_X1 U541 ( .A(n606), .B(n530), .ZN(n405) );
  AND2_X1 U542 ( .A1(n384), .A2(n383), .ZN(n382) );
  NAND2_X1 U543 ( .A1(n406), .A2(n414), .ZN(n411) );
  NAND2_X1 U544 ( .A1(n357), .A2(n388), .ZN(n476) );
  XNOR2_X1 U545 ( .A(n590), .B(n362), .ZN(n377) );
  XNOR2_X2 U546 ( .A(n563), .B(n562), .ZN(n749) );
  INV_X1 U547 ( .A(n570), .ZN(n517) );
  NAND2_X1 U548 ( .A1(n379), .A2(n407), .ZN(n413) );
  NAND2_X1 U549 ( .A1(n464), .A2(n380), .ZN(n388) );
  NOR2_X1 U550 ( .A1(n663), .A2(n387), .ZN(n380) );
  OR2_X1 U551 ( .A1(n575), .A2(n381), .ZN(n385) );
  NAND2_X1 U552 ( .A1(n663), .A2(n386), .ZN(n384) );
  NAND2_X1 U553 ( .A1(n748), .A2(n398), .ZN(n392) );
  AND2_X1 U554 ( .A1(n610), .A2(n395), .ZN(n394) );
  NAND2_X1 U555 ( .A1(n752), .A2(KEYINPUT46), .ZN(n395) );
  NOR2_X1 U556 ( .A1(n752), .A2(KEYINPUT46), .ZN(n397) );
  INV_X1 U557 ( .A(KEYINPUT46), .ZN(n398) );
  NOR2_X1 U558 ( .A1(n465), .A2(n721), .ZN(G54) );
  XNOR2_X2 U559 ( .A(n399), .B(G472), .ZN(n597) );
  NAND2_X1 U560 ( .A1(n401), .A2(n729), .ZN(n730) );
  XNOR2_X1 U561 ( .A(n402), .B(G134), .ZN(n489) );
  NOR2_X2 U562 ( .A1(n405), .A2(n537), .ZN(n538) );
  NOR2_X1 U563 ( .A1(n611), .A2(n405), .ZN(n656) );
  INV_X1 U564 ( .A(n415), .ZN(n406) );
  NAND2_X1 U565 ( .A1(n412), .A2(n363), .ZN(n410) );
  AND2_X1 U566 ( .A1(n415), .A2(KEYINPUT80), .ZN(n409) );
  XNOR2_X1 U567 ( .A(n416), .B(n506), .ZN(n507) );
  NOR2_X2 U568 ( .A1(n447), .A2(n451), .ZN(n562) );
  XNOR2_X2 U569 ( .A(n417), .B(G146), .ZN(n523) );
  XNOR2_X2 U570 ( .A(n571), .B(KEYINPUT31), .ZN(n663) );
  NOR2_X1 U571 ( .A1(n425), .A2(n606), .ZN(n608) );
  NOR2_X2 U572 ( .A1(n403), .A2(n609), .ZN(n665) );
  NOR2_X2 U573 ( .A1(n454), .A2(n455), .ZN(n631) );
  XNOR2_X2 U574 ( .A(n445), .B(n444), .ZN(n454) );
  INV_X1 U575 ( .A(n567), .ZN(n652) );
  NAND2_X1 U576 ( .A1(n630), .A2(n629), .ZN(n455) );
  XNOR2_X1 U577 ( .A(n618), .B(KEYINPUT70), .ZN(n429) );
  XNOR2_X1 U578 ( .A(n430), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U579 ( .A1(n710), .A2(n721), .ZN(n430) );
  XNOR2_X1 U580 ( .A(n432), .B(n643), .ZN(G57) );
  XNOR2_X1 U581 ( .A(n433), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U582 ( .A1(n717), .A2(n721), .ZN(n433) );
  INV_X1 U583 ( .A(n577), .ZN(n579) );
  NOR2_X1 U584 ( .A1(n662), .A2(n660), .ZN(n580) );
  NAND2_X1 U585 ( .A1(n436), .A2(n434), .ZN(n617) );
  NAND2_X1 U586 ( .A1(n656), .A2(n463), .ZN(n435) );
  XNOR2_X1 U587 ( .A(n438), .B(n437), .ZN(n436) );
  INV_X1 U588 ( .A(KEYINPUT71), .ZN(n437) );
  NAND2_X1 U589 ( .A1(n439), .A2(n656), .ZN(n438) );
  XNOR2_X1 U590 ( .A(n612), .B(KEYINPUT72), .ZN(n439) );
  XNOR2_X1 U591 ( .A(n557), .B(n558), .ZN(n443) );
  INV_X1 U592 ( .A(n454), .ZN(n723) );
  NAND2_X1 U593 ( .A1(n449), .A2(n353), .ZN(n447) );
  NAND2_X1 U594 ( .A1(n682), .A2(n450), .ZN(n449) );
  NOR2_X1 U595 ( .A1(n682), .A2(n360), .ZN(n451) );
  XNOR2_X1 U596 ( .A(n455), .B(n737), .ZN(n738) );
  NAND2_X1 U597 ( .A1(n354), .A2(G469), .ZN(n467) );
  NAND2_X1 U598 ( .A1(n354), .A2(G478), .ZN(n718) );
  NAND2_X1 U599 ( .A1(n613), .A2(n684), .ZN(n593) );
  INV_X1 U600 ( .A(n464), .ZN(n645) );
  XNOR2_X1 U601 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X2 U602 ( .A1(n707), .A2(n526), .ZN(n528) );
  XNOR2_X1 U603 ( .A(KEYINPUT59), .B(KEYINPUT83), .ZN(n474) );
  NOR2_X1 U604 ( .A1(n603), .A2(n347), .ZN(n475) );
  INV_X1 U605 ( .A(n668), .ZN(n628) );
  INV_X1 U606 ( .A(KEYINPUT87), .ZN(n539) );
  NOR2_X1 U607 ( .A1(n753), .A2(n628), .ZN(n629) );
  INV_X1 U608 ( .A(KEYINPUT36), .ZN(n607) );
  XNOR2_X1 U609 ( .A(n716), .B(n715), .ZN(n717) );
  INV_X1 U610 ( .A(KEYINPUT119), .ZN(n636) );
  XOR2_X1 U611 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n478) );
  XNOR2_X1 U612 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U613 ( .A(n736), .B(n481), .Z(n484) );
  NAND2_X1 U614 ( .A1(G234), .A2(n722), .ZN(n482) );
  XOR2_X1 U615 ( .A(KEYINPUT8), .B(n482), .Z(n546) );
  NAND2_X1 U616 ( .A1(G221), .A2(n546), .ZN(n483) );
  XOR2_X1 U617 ( .A(n484), .B(n483), .Z(n634) );
  INV_X1 U618 ( .A(KEYINPUT35), .ZN(n563) );
  XNOR2_X2 U619 ( .A(n485), .B(G143), .ZN(n543) );
  XNOR2_X1 U620 ( .A(n487), .B(KEYINPUT66), .ZN(n550) );
  INV_X1 U621 ( .A(n550), .ZN(n488) );
  XNOR2_X1 U622 ( .A(n490), .B(G104), .ZN(n493) );
  AND2_X1 U623 ( .A1(G227), .A2(n722), .ZN(n494) );
  XNOR2_X1 U624 ( .A(n520), .B(n494), .ZN(n495) );
  XOR2_X1 U625 ( .A(KEYINPUT76), .B(KEYINPUT88), .Z(n496) );
  INV_X1 U626 ( .A(G469), .ZN(n497) );
  NOR2_X1 U627 ( .A1(n634), .A2(G902), .ZN(n503) );
  XOR2_X1 U628 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n501) );
  INV_X1 U629 ( .A(n526), .ZN(n632) );
  NAND2_X1 U630 ( .A1(G234), .A2(n632), .ZN(n499) );
  XNOR2_X1 U631 ( .A(KEYINPUT20), .B(n499), .ZN(n504) );
  NAND2_X1 U632 ( .A1(n504), .A2(G217), .ZN(n500) );
  XNOR2_X1 U633 ( .A(n501), .B(n500), .ZN(n502) );
  NAND2_X1 U634 ( .A1(n504), .A2(G221), .ZN(n505) );
  XOR2_X1 U635 ( .A(KEYINPUT21), .B(n505), .Z(n669) );
  INV_X1 U636 ( .A(n669), .ZN(n564) );
  NOR2_X1 U637 ( .A1(n592), .A2(n564), .ZN(n673) );
  XNOR2_X1 U638 ( .A(n510), .B(n509), .ZN(n514) );
  NAND2_X1 U639 ( .A1(n552), .A2(G210), .ZN(n511) );
  XNOR2_X1 U640 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U641 ( .A(n514), .B(n513), .Z(n515) );
  NAND2_X1 U642 ( .A1(n517), .A2(n603), .ZN(n518) );
  XOR2_X1 U643 ( .A(G116), .B(G107), .Z(n542) );
  NAND2_X1 U644 ( .A1(G224), .A2(n722), .ZN(n525) );
  NAND2_X1 U645 ( .A1(G210), .A2(n529), .ZN(n527) );
  XNOR2_X2 U646 ( .A(n528), .B(n527), .ZN(n625) );
  NAND2_X1 U647 ( .A1(G214), .A2(n529), .ZN(n683) );
  NAND2_X1 U648 ( .A1(n625), .A2(n683), .ZN(n606) );
  NAND2_X1 U649 ( .A1(G237), .A2(G234), .ZN(n531) );
  XNOR2_X1 U650 ( .A(n531), .B(KEYINPUT14), .ZN(n534) );
  NAND2_X1 U651 ( .A1(G952), .A2(n534), .ZN(n698) );
  NOR2_X1 U652 ( .A1(n698), .A2(G953), .ZN(n532) );
  XNOR2_X1 U653 ( .A(n532), .B(KEYINPUT85), .ZN(n587) );
  INV_X1 U654 ( .A(n587), .ZN(n536) );
  NOR2_X1 U655 ( .A1(G898), .A2(n722), .ZN(n533) );
  XOR2_X1 U656 ( .A(KEYINPUT86), .B(n533), .Z(n729) );
  NAND2_X1 U657 ( .A1(G902), .A2(n534), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n729), .A2(n585), .ZN(n535) );
  NOR2_X1 U659 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U660 ( .A(n541), .B(n540), .ZN(n545) );
  XNOR2_X1 U661 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U662 ( .A1(G217), .A2(n546), .ZN(n547) );
  XNOR2_X1 U663 ( .A(n548), .B(n547), .ZN(n719) );
  NOR2_X1 U664 ( .A1(G902), .A2(n719), .ZN(n549) );
  XNOR2_X1 U665 ( .A(G478), .B(n549), .ZN(n576) );
  INV_X1 U666 ( .A(n576), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n551), .B(n550), .ZN(n557) );
  XOR2_X1 U668 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n554) );
  NAND2_X1 U669 ( .A1(n552), .A2(G214), .ZN(n553) );
  XNOR2_X1 U670 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U671 ( .A1(G902), .A2(n714), .ZN(n560) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(G475), .ZN(n559) );
  NAND2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n561) );
  XNOR2_X1 U674 ( .A(n561), .B(KEYINPUT101), .ZN(n615) );
  NAND2_X1 U675 ( .A1(n579), .A2(n576), .ZN(n687) );
  NOR2_X1 U676 ( .A1(n687), .A2(n564), .ZN(n565) );
  NOR2_X1 U677 ( .A1(n603), .A2(n568), .ZN(n569) );
  NAND2_X1 U678 ( .A1(n347), .A2(n569), .ZN(n644) );
  INV_X1 U679 ( .A(n597), .ZN(n672) );
  INV_X1 U680 ( .A(n601), .ZN(n591) );
  AND2_X1 U681 ( .A1(n673), .A2(n601), .ZN(n572) );
  XNOR2_X1 U682 ( .A(n574), .B(KEYINPUT91), .ZN(n575) );
  NOR2_X1 U683 ( .A1(n577), .A2(n576), .ZN(n662) );
  NOR2_X1 U684 ( .A1(n749), .A2(KEYINPUT44), .ZN(n581) );
  XNOR2_X1 U685 ( .A(n582), .B(KEYINPUT81), .ZN(n583) );
  NOR2_X1 U686 ( .A1(G900), .A2(n585), .ZN(n586) );
  NAND2_X1 U687 ( .A1(G953), .A2(n586), .ZN(n588) );
  NAND2_X1 U688 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U689 ( .A1(n589), .A2(n669), .ZN(n595) );
  NAND2_X1 U690 ( .A1(n597), .A2(n683), .ZN(n590) );
  NAND2_X1 U691 ( .A1(n684), .A2(n683), .ZN(n688) );
  XNOR2_X1 U692 ( .A(KEYINPUT41), .B(n594), .ZN(n699) );
  XNOR2_X1 U693 ( .A(KEYINPUT68), .B(n595), .ZN(n596) );
  XNOR2_X1 U694 ( .A(KEYINPUT28), .B(KEYINPUT104), .ZN(n598) );
  NOR2_X1 U695 ( .A1(n699), .A2(n611), .ZN(n602) );
  AND2_X1 U696 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U697 ( .A1(n660), .A2(n605), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(n665), .ZN(n610) );
  NOR2_X1 U700 ( .A1(KEYINPUT47), .A2(n689), .ZN(n612) );
  AND2_X1 U701 ( .A1(n431), .A2(n613), .ZN(n614) );
  NAND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U703 ( .A(KEYINPUT103), .B(n616), .ZN(n750) );
  XNOR2_X1 U704 ( .A(n619), .B(KEYINPUT48), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n620), .A2(n662), .ZN(n621) );
  XOR2_X1 U706 ( .A(KEYINPUT106), .B(n621), .Z(n753) );
  NOR2_X1 U707 ( .A1(n674), .A2(n622), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n623), .A2(n683), .ZN(n624) );
  XNOR2_X1 U709 ( .A(n624), .B(KEYINPUT43), .ZN(n627) );
  INV_X1 U710 ( .A(n431), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n668) );
  XNOR2_X1 U712 ( .A(n633), .B(n634), .ZN(n635) );
  NOR2_X2 U713 ( .A1(n635), .A2(n721), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(n636), .ZN(G66) );
  XOR2_X1 U715 ( .A(KEYINPUT62), .B(KEYINPUT107), .Z(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT63), .B(KEYINPUT108), .Z(n643) );
  XNOR2_X1 U717 ( .A(G101), .B(n644), .ZN(G3) );
  XOR2_X1 U718 ( .A(G104), .B(KEYINPUT109), .Z(n647) );
  NAND2_X1 U719 ( .A1(n645), .A2(n660), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G6) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT27), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n649) );
  NAND2_X1 U723 ( .A1(n645), .A2(n662), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(G9) );
  XOR2_X1 U726 ( .A(n652), .B(G110), .Z(G12) );
  XOR2_X1 U727 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n654) );
  NAND2_X1 U728 ( .A1(n656), .A2(n662), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(n655) );
  XOR2_X1 U730 ( .A(G128), .B(n655), .Z(G30) );
  XOR2_X1 U731 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n658) );
  NAND2_X1 U732 ( .A1(n656), .A2(n660), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U734 ( .A(G146), .B(n659), .ZN(G48) );
  NAND2_X1 U735 ( .A1(n663), .A2(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(G113), .ZN(G15) );
  NAND2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(G116), .ZN(G18) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT37), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n666), .B(KEYINPUT114), .ZN(n667) );
  XNOR2_X1 U741 ( .A(G125), .B(n667), .ZN(G27) );
  XNOR2_X1 U742 ( .A(G140), .B(n668), .ZN(G42) );
  XOR2_X1 U743 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n696) );
  NOR2_X1 U744 ( .A1(n347), .A2(n669), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(KEYINPUT49), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U751 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NOR2_X1 U752 ( .A1(n699), .A2(n681), .ZN(n694) );
  INV_X1 U753 ( .A(n682), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U755 ( .A(KEYINPUT115), .B(n685), .Z(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n700), .A2(n692), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U761 ( .A(n696), .B(n695), .Z(n697) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U766 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n706) );
  XNOR2_X1 U767 ( .A(n707), .B(n706), .ZN(n708) );
  XOR2_X1 U768 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n713) );
  XNOR2_X1 U769 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n721), .A2(n720), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(KEYINPUT120), .ZN(n728) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n725), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G898), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n731) );
  XOR2_X1 U778 ( .A(n731), .B(n730), .Z(G69) );
  XNOR2_X1 U779 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n734) );
  XNOR2_X1 U780 ( .A(n732), .B(KEYINPUT88), .ZN(n733) );
  XNOR2_X1 U781 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n736), .B(n735), .ZN(n741) );
  INV_X1 U783 ( .A(n741), .ZN(n737) );
  NOR2_X1 U784 ( .A1(G953), .A2(n738), .ZN(n739) );
  XNOR2_X1 U785 ( .A(KEYINPUT123), .B(n739), .ZN(n746) );
  XNOR2_X1 U786 ( .A(G227), .B(KEYINPUT124), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(G953), .ZN(n744) );
  XOR2_X1 U790 ( .A(KEYINPUT125), .B(n744), .Z(n745) );
  NAND2_X1 U791 ( .A1(n746), .A2(n745), .ZN(G72) );
  XOR2_X1 U792 ( .A(G131), .B(KEYINPUT126), .Z(n747) );
  XNOR2_X1 U793 ( .A(n748), .B(n747), .ZN(G33) );
  XOR2_X1 U794 ( .A(n749), .B(G122), .Z(G24) );
  XOR2_X1 U795 ( .A(G143), .B(n750), .Z(G45) );
  XOR2_X1 U796 ( .A(n751), .B(G119), .Z(G21) );
  XOR2_X1 U797 ( .A(G137), .B(n752), .Z(G39) );
  XOR2_X1 U798 ( .A(G134), .B(n753), .Z(G36) );
endmodule

