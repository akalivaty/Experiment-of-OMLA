

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(G2105), .A2(n516), .ZN(n874) );
  INV_X1 U552 ( .A(KEYINPUT23), .ZN(n533) );
  NOR2_X1 U553 ( .A1(n989), .A2(n682), .ZN(n684) );
  AND2_X1 U554 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U555 ( .A1(n539), .A2(n538), .ZN(G160) );
  INV_X1 U556 ( .A(KEYINPUT64), .ZN(n683) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n700) );
  NOR2_X1 U558 ( .A1(n718), .A2(n717), .ZN(n719) );
  BUF_X1 U559 ( .A(n679), .Z(n732) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n722) );
  NOR2_X1 U561 ( .A1(G1966), .A2(n762), .ZN(n724) );
  NOR2_X1 U562 ( .A1(n676), .A2(n768), .ZN(n706) );
  INV_X1 U563 ( .A(n970), .ZN(n752) );
  NOR2_X1 U564 ( .A1(n751), .A2(n752), .ZN(n753) );
  XNOR2_X1 U565 ( .A(G2104), .B(KEYINPUT66), .ZN(n524) );
  NOR2_X1 U566 ( .A1(n525), .A2(G2105), .ZN(n532) );
  BUF_X1 U567 ( .A(n532), .Z(n870) );
  XNOR2_X1 U568 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U569 ( .A(KEYINPUT65), .B(n540), .Z(n649) );
  NAND2_X1 U570 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U571 ( .A1(n528), .A2(n527), .ZN(G164) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U573 ( .A1(G114), .A2(n876), .ZN(n518) );
  XOR2_X1 U574 ( .A(G2104), .B(KEYINPUT66), .Z(n516) );
  NAND2_X1 U575 ( .A1(G126), .A2(n874), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U577 ( .A(n519), .B(KEYINPUT83), .ZN(n523) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X1 U579 ( .A(KEYINPUT17), .B(n520), .Z(n521) );
  XNOR2_X1 U580 ( .A(KEYINPUT68), .B(n521), .ZN(n529) );
  NAND2_X1 U581 ( .A1(G138), .A2(n529), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n523), .A2(n522), .ZN(n528) );
  INV_X1 U583 ( .A(n524), .ZN(n525) );
  NAND2_X1 U584 ( .A1(G102), .A2(n870), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT84), .B(n526), .Z(n527) );
  NAND2_X1 U586 ( .A1(G113), .A2(n876), .ZN(n531) );
  BUF_X1 U587 ( .A(n529), .Z(n871) );
  NAND2_X1 U588 ( .A1(G137), .A2(n871), .ZN(n530) );
  AND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n532), .A2(G101), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n874), .A2(G125), .ZN(n535) );
  XNOR2_X1 U592 ( .A(KEYINPUT67), .B(n537), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n622) );
  NOR2_X1 U594 ( .A1(G651), .A2(n622), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n649), .A2(G52), .ZN(n541) );
  XOR2_X1 U596 ( .A(KEYINPUT71), .B(n541), .Z(n544) );
  INV_X1 U597 ( .A(G651), .ZN(n547) );
  NOR2_X1 U598 ( .A1(G543), .A2(n547), .ZN(n542) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n542), .Z(n643) );
  NAND2_X1 U600 ( .A1(n643), .A2(G64), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT72), .B(n545), .ZN(n552) );
  NOR2_X1 U603 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U604 ( .A1(n642), .A2(G90), .ZN(n546) );
  XOR2_X1 U605 ( .A(KEYINPUT73), .B(n546), .Z(n549) );
  NOR2_X1 U606 ( .A1(n622), .A2(n547), .ZN(n640) );
  NAND2_X1 U607 ( .A1(n640), .A2(G77), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U610 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U611 ( .A1(G111), .A2(n876), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G135), .A2(n871), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n874), .A2(G123), .ZN(n555) );
  XOR2_X1 U615 ( .A(KEYINPUT18), .B(n555), .Z(n556) );
  NOR2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n870), .A2(G99), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n912) );
  XNOR2_X1 U619 ( .A(G2096), .B(n912), .ZN(n560) );
  OR2_X1 U620 ( .A1(G2100), .A2(n560), .ZN(G156) );
  NAND2_X1 U621 ( .A1(G91), .A2(n642), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G65), .A2(n643), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G78), .A2(n640), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G53), .A2(n649), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n978) );
  INV_X1 U628 ( .A(n978), .ZN(G299) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(n649), .A2(G51), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT78), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G63), .A2(n643), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT6), .B(n570), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n642), .A2(G89), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G76), .A2(n640), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT77), .B(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT5), .B(n575), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT7), .B(n578), .Z(G168) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G94), .A2(G452), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT74), .B(n579), .Z(G173) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n580) );
  XOR2_X1 U649 ( .A(n580), .B(KEYINPUT10), .Z(n820) );
  NAND2_X1 U650 ( .A1(n820), .A2(G567), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n581), .B(KEYINPUT11), .ZN(n582) );
  XNOR2_X1 U652 ( .A(KEYINPUT75), .B(n582), .ZN(G234) );
  NAND2_X1 U653 ( .A1(G56), .A2(n643), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U655 ( .A1(n642), .A2(G81), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G68), .A2(n640), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n649), .A2(G43), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n989) );
  INV_X1 U663 ( .A(G860), .ZN(n611) );
  OR2_X1 U664 ( .A1(n989), .A2(n611), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  INV_X1 U666 ( .A(G868), .ZN(n602) );
  NOR2_X1 U667 ( .A1(G301), .A2(n602), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G92), .A2(n642), .ZN(n593) );
  NAND2_X1 U669 ( .A1(G66), .A2(n643), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G79), .A2(n640), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G54), .A2(n649), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT15), .B(n598), .Z(n599) );
  XOR2_X1 U676 ( .A(KEYINPUT76), .B(n599), .Z(n975) );
  NOR2_X1 U677 ( .A1(n975), .A2(G868), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(G284) );
  NOR2_X1 U679 ( .A1(G286), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n611), .A2(G559), .ZN(n605) );
  INV_X1 U683 ( .A(n975), .ZN(n891) );
  NAND2_X1 U684 ( .A1(n605), .A2(n891), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n989), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n891), .A2(G868), .ZN(n607) );
  NOR2_X1 U688 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U689 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U690 ( .A1(n891), .A2(G559), .ZN(n610) );
  XOR2_X1 U691 ( .A(n989), .B(n610), .Z(n657) );
  NAND2_X1 U692 ( .A1(n611), .A2(n657), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G93), .A2(n642), .ZN(n613) );
  NAND2_X1 U694 ( .A1(G67), .A2(n643), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G80), .A2(n640), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G55), .A2(n649), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n659) );
  XOR2_X1 U700 ( .A(n618), .B(n659), .Z(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n649), .ZN(n620) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n643), .A2(n621), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n622), .A2(G87), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G85), .A2(n642), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G72), .A2(n640), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U710 ( .A(KEYINPUT69), .B(n627), .Z(n630) );
  NAND2_X1 U711 ( .A1(G60), .A2(n643), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT70), .B(n628), .Z(n629) );
  NOR2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n649), .A2(G47), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U716 ( .A1(G88), .A2(n642), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G75), .A2(n640), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U719 ( .A(KEYINPUT80), .B(n635), .Z(n639) );
  NAND2_X1 U720 ( .A1(G62), .A2(n643), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G50), .A2(n649), .ZN(n636) );
  AND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(G303) );
  INV_X1 U724 ( .A(G303), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G73), .A2(n640), .ZN(n641) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n641), .Z(n648) );
  NAND2_X1 U727 ( .A1(G86), .A2(n642), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G61), .A2(n643), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U730 ( .A(KEYINPUT79), .B(n646), .Z(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n649), .A2(G48), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(G305) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XOR2_X1 U735 ( .A(G299), .B(n659), .Z(n654) );
  XOR2_X1 U736 ( .A(G290), .B(G166), .Z(n652) );
  XNOR2_X1 U737 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U738 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n656), .B(n655), .ZN(n889) );
  XNOR2_X1 U740 ( .A(n657), .B(n889), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n658), .A2(G868), .ZN(n661) );
  OR2_X1 U742 ( .A1(G868), .A2(n659), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n663), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n664) );
  XNOR2_X1 U748 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U749 ( .A1(G2072), .A2(n666), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U752 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U753 ( .A1(G108), .A2(n668), .ZN(n825) );
  NAND2_X1 U754 ( .A1(n825), .A2(G567), .ZN(n674) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n669) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n670), .A2(G96), .ZN(n671) );
  NOR2_X1 U758 ( .A1(G218), .A2(n671), .ZN(n672) );
  XOR2_X1 U759 ( .A(KEYINPUT82), .B(n672), .Z(n826) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n826), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n827) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U763 ( .A1(n827), .A2(n675), .ZN(n824) );
  NAND2_X1 U764 ( .A1(n824), .A2(G36), .ZN(G176) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n767) );
  INV_X1 U766 ( .A(n767), .ZN(n676) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U768 ( .A(n706), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G8), .A2(n679), .ZN(n762) );
  XNOR2_X1 U770 ( .A(G1996), .B(KEYINPUT93), .ZN(n945) );
  NOR2_X1 U771 ( .A1(n679), .A2(n945), .ZN(n678) );
  XOR2_X1 U772 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n677) );
  XNOR2_X1 U773 ( .A(n678), .B(n677), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n732), .A2(G1341), .ZN(n680) );
  NAND2_X1 U775 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U776 ( .A(n684), .B(n683), .ZN(n688) );
  XNOR2_X1 U777 ( .A(n706), .B(KEYINPUT91), .ZN(n694) );
  INV_X1 U778 ( .A(n694), .ZN(n708) );
  NAND2_X1 U779 ( .A1(G2067), .A2(n708), .ZN(n686) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n732), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n686), .A2(n685), .ZN(n689) );
  OR2_X1 U782 ( .A1(n689), .A2(n975), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n975), .A2(n689), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n698) );
  INV_X1 U786 ( .A(G2072), .ZN(n930) );
  NOR2_X1 U787 ( .A1(n694), .A2(n930), .ZN(n693) );
  XNOR2_X1 U788 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U789 ( .A(n693), .B(n692), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n694), .A2(G1956), .ZN(n695) );
  AND2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n978), .A2(n699), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n699), .A2(n978), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U798 ( .A(n705), .B(n704), .ZN(n712) );
  NOR2_X1 U799 ( .A1(n706), .A2(G1961), .ZN(n707) );
  XOR2_X1 U800 ( .A(KEYINPUT90), .B(n707), .Z(n710) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U802 ( .A1(n708), .A2(n944), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n716), .A2(G171), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n721) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n732), .ZN(n725) );
  NOR2_X1 U807 ( .A1(n724), .A2(n725), .ZN(n713) );
  NAND2_X1 U808 ( .A1(G8), .A2(n713), .ZN(n714) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U810 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U811 ( .A1(G171), .A2(n716), .ZN(n717) );
  XOR2_X1 U812 ( .A(KEYINPUT31), .B(n719), .Z(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n730) );
  XNOR2_X1 U814 ( .A(n730), .B(n722), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U816 ( .A1(n725), .A2(G8), .ZN(n726) );
  XOR2_X1 U817 ( .A(KEYINPUT89), .B(n726), .Z(n727) );
  NAND2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n743) );
  AND2_X1 U819 ( .A1(G286), .A2(G8), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n740) );
  INV_X1 U821 ( .A(G8), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n762), .ZN(n731) );
  XOR2_X1 U823 ( .A(KEYINPUT97), .B(n731), .Z(n734) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U826 ( .A(n735), .B(KEYINPUT98), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n741), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n749), .A2(n744), .ZN(n972) );
  NAND2_X1 U834 ( .A1(n758), .A2(n972), .ZN(n745) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NAND2_X1 U836 ( .A1(n745), .A2(n977), .ZN(n746) );
  NOR2_X1 U837 ( .A1(n762), .A2(n746), .ZN(n747) );
  NOR2_X1 U838 ( .A1(KEYINPUT33), .A2(n747), .ZN(n748) );
  XNOR2_X1 U839 ( .A(n748), .B(KEYINPUT99), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n762), .A2(n750), .ZN(n751) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n970) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT100), .ZN(n766) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U846 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U848 ( .A1(n759), .A2(n762), .ZN(n764) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U850 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  NOR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n802) );
  BUF_X1 U854 ( .A(n767), .Z(n769) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n813) );
  XNOR2_X1 U856 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U857 ( .A1(G104), .A2(n870), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G140), .A2(n871), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n772), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G116), .A2(n876), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G128), .A2(n874), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U864 ( .A(KEYINPUT85), .B(n775), .ZN(n776) );
  XNOR2_X1 U865 ( .A(KEYINPUT35), .B(n776), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n779), .ZN(n886) );
  NOR2_X1 U868 ( .A1(n810), .A2(n886), .ZN(n925) );
  NAND2_X1 U869 ( .A1(n813), .A2(n925), .ZN(n808) );
  NAND2_X1 U870 ( .A1(G107), .A2(n876), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G131), .A2(n871), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n870), .A2(G95), .ZN(n782) );
  XOR2_X1 U874 ( .A(KEYINPUT86), .B(n782), .Z(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n874), .A2(G119), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n883) );
  AND2_X1 U878 ( .A1(n883), .A2(G1991), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G117), .A2(n876), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G141), .A2(n871), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G105), .A2(n870), .ZN(n789) );
  XNOR2_X1 U883 ( .A(n789), .B(KEYINPUT38), .ZN(n790) );
  XNOR2_X1 U884 ( .A(n790), .B(KEYINPUT87), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n874), .A2(G129), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n865) );
  AND2_X1 U888 ( .A1(n865), .A2(G1996), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n913) );
  XOR2_X1 U890 ( .A(n813), .B(KEYINPUT88), .Z(n797) );
  NOR2_X1 U891 ( .A1(n913), .A2(n797), .ZN(n805) );
  INV_X1 U892 ( .A(n805), .ZN(n798) );
  AND2_X1 U893 ( .A1(n808), .A2(n798), .ZN(n800) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U895 ( .A1(n973), .A2(n813), .ZN(n799) );
  AND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n816) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n865), .ZN(n917) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n883), .ZN(n915) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n915), .A2(n803), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n917), .A2(n806), .ZN(n807) );
  XNOR2_X1 U904 ( .A(KEYINPUT39), .B(n807), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n812) );
  AND2_X1 U906 ( .A1(n886), .A2(n810), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT101), .ZN(n927) );
  NAND2_X1 U908 ( .A1(n812), .A2(n927), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n819) );
  XOR2_X1 U911 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT102), .B(n817), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n819), .B(n818), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n820), .ZN(G217) );
  INV_X1 U915 ( .A(n820), .ZN(G223) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n821) );
  XOR2_X1 U917 ( .A(KEYINPUT106), .B(n821), .Z(n822) );
  NAND2_X1 U918 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n827), .ZN(G319) );
  XOR2_X1 U928 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n829) );
  XNOR2_X1 U929 ( .A(KEYINPUT108), .B(G2678), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2090), .Z(n831) );
  XOR2_X1 U932 ( .A(G2067), .B(n930), .Z(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U934 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U935 ( .A(G2096), .B(G2100), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U937 ( .A(G2084), .B(G2078), .Z(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1981), .B(G1961), .Z(n839) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1956), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n840), .B(G2474), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1976), .Z(n844) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1971), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G112), .A2(n876), .ZN(n848) );
  NAND2_X1 U950 ( .A1(G136), .A2(n871), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n874), .A2(G124), .ZN(n849) );
  XNOR2_X1 U953 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U954 ( .A1(G100), .A2(n870), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U956 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U957 ( .A1(G118), .A2(n876), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G130), .A2(n874), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G106), .A2(n870), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G142), .A2(n871), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U963 ( .A(n858), .B(KEYINPUT45), .Z(n859) );
  NOR2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(n861), .Z(n862) );
  XNOR2_X1 U966 ( .A(KEYINPUT112), .B(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n912), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n868) );
  XNOR2_X1 U970 ( .A(G164), .B(G160), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(n869), .B(G162), .Z(n885) );
  NAND2_X1 U973 ( .A1(G103), .A2(n870), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G139), .A2(n871), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n882) );
  NAND2_X1 U976 ( .A1(n874), .A2(G127), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(KEYINPUT110), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G115), .A2(n876), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(KEYINPUT47), .B(n879), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n880), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n929) );
  XOR2_X1 U983 ( .A(n883), .B(n929), .Z(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U986 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U987 ( .A(G301), .B(G286), .Z(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n989), .B(n891), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U991 ( .A1(G37), .A2(n894), .ZN(G397) );
  XNOR2_X1 U992 ( .A(G2427), .B(KEYINPUT104), .ZN(n904) );
  XOR2_X1 U993 ( .A(G2430), .B(G2446), .Z(n896) );
  XNOR2_X1 U994 ( .A(G2435), .B(G2438), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U996 ( .A(G2454), .B(KEYINPUT105), .Z(n898) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U999 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G2451), .B(G2443), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n905), .A2(G14), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(n911), .ZN(G401) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n923) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n921) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1018 ( .A(KEYINPUT113), .B(n918), .Z(n919) );
  XNOR2_X1 U1019 ( .A(KEYINPUT51), .B(n919), .ZN(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n926), .B(KEYINPUT114), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n936) );
  XOR2_X1 U1025 ( .A(n930), .B(n929), .Z(n932) );
  XNOR2_X1 U1026 ( .A(G164), .B(G2078), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1028 ( .A(KEYINPUT115), .B(n933), .Z(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n934), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1035 ( .A(G2084), .B(G34), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(KEYINPUT54), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n962) );
  XNOR2_X1 U1039 ( .A(G27), .B(n944), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(n945), .B(G32), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G33), .B(KEYINPUT118), .ZN(n946) );
  XOR2_X1 U1042 ( .A(n946), .B(G2072), .Z(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1044 ( .A(KEYINPUT117), .B(G2067), .Z(n949) );
  XNOR2_X1 U1045 ( .A(G26), .B(n949), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT119), .B(n954), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G25), .B(G1991), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(KEYINPUT116), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(n959), .B(KEYINPUT120), .Z(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1056 ( .A(KEYINPUT55), .B(n963), .Z(n965) );
  INV_X1 U1057 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n966), .ZN(n1024) );
  XNOR2_X1 U1060 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n967) );
  XOR2_X1 U1061 ( .A(G16), .B(n967), .Z(n996) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G168), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT122), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT57), .B(n971), .ZN(n994) );
  INV_X1 U1066 ( .A(n972), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n986) );
  XOR2_X1 U1068 ( .A(G1348), .B(n975), .Z(n982) );
  NAND2_X1 U1069 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n980) );
  XOR2_X1 U1071 ( .A(G1956), .B(n978), .Z(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G1961), .B(G171), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(KEYINPUT123), .B(n987), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G1341), .B(KEYINPUT124), .Z(n988) );
  XNOR2_X1 U1079 ( .A(n989), .B(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n992), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1022) );
  INV_X1 U1084 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1085 ( .A(G1976), .B(G23), .Z(n998) );
  XOR2_X1 U1086 ( .A(G1971), .B(G22), .Z(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G24), .B(G1986), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT58), .B(n1001), .Z(n1017) );
  XOR2_X1 U1091 ( .A(G1966), .B(G21), .Z(n1011) );
  XNOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(G1961), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(G5), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .ZN(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

