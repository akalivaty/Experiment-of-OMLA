

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782;

  AND2_X1 U374 ( .A1(n593), .A2(n409), .ZN(n408) );
  XNOR2_X1 U375 ( .A(n463), .B(G104), .ZN(n531) );
  XNOR2_X1 U376 ( .A(n387), .B(n364), .ZN(n386) );
  NAND2_X1 U377 ( .A1(n386), .A2(n657), .ZN(n768) );
  XNOR2_X1 U378 ( .A(n465), .B(n464), .ZN(n545) );
  XOR2_X1 U379 ( .A(KEYINPUT89), .B(KEYINPUT78), .Z(n352) );
  INV_X2 U380 ( .A(n681), .ZN(n752) );
  INV_X1 U381 ( .A(n576), .ZN(n438) );
  NAND2_X2 U382 ( .A1(n456), .A2(n363), .ZN(n427) );
  NAND2_X1 U383 ( .A1(n702), .A2(n700), .ZN(n391) );
  NOR2_X2 U384 ( .A1(n722), .A2(n721), .ZN(n585) );
  XNOR2_X2 U385 ( .A(G119), .B(G116), .ZN(n453) );
  NAND2_X1 U386 ( .A1(n410), .A2(n408), .ZN(n407) );
  NOR2_X1 U387 ( .A1(n433), .A2(n779), .ZN(n388) );
  NOR2_X1 U388 ( .A1(n646), .A2(n618), .ZN(n619) );
  AND2_X1 U389 ( .A1(n400), .A2(n397), .ZN(n396) );
  NOR2_X1 U390 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U391 ( .A(n414), .B(KEYINPUT105), .ZN(n634) );
  XNOR2_X1 U392 ( .A(n612), .B(KEYINPUT1), .ZN(n722) );
  OR2_X2 U393 ( .A1(n583), .A2(n584), .ZN(n700) );
  XNOR2_X1 U394 ( .A(n559), .B(n449), .ZN(n725) );
  XNOR2_X1 U395 ( .A(n458), .B(n496), .ZN(n584) );
  NAND2_X2 U396 ( .A1(n379), .A2(n376), .ZN(n612) );
  XNOR2_X1 U397 ( .A(n546), .B(n680), .ZN(n610) );
  AND2_X1 U398 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U399 ( .A(n667), .B(n666), .ZN(n668) );
  OR2_X1 U400 ( .A1(n754), .A2(n377), .ZN(n376) );
  NAND2_X1 U401 ( .A1(n535), .A2(n378), .ZN(n377) );
  XNOR2_X1 U402 ( .A(G113), .B(KEYINPUT3), .ZN(n452) );
  INV_X1 U403 ( .A(G953), .ZN(n527) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(G902), .ZN(n659) );
  BUF_X2 U405 ( .A(n633), .Z(n654) );
  XNOR2_X1 U406 ( .A(n367), .B(n366), .ZN(n519) );
  INV_X1 U407 ( .A(KEYINPUT92), .ZN(n366) );
  NAND2_X1 U408 ( .A1(n450), .A2(n448), .ZN(n620) );
  NOR2_X1 U409 ( .A1(n629), .A2(n451), .ZN(n450) );
  NOR2_X1 U410 ( .A1(n584), .A2(n582), .ZN(n414) );
  INV_X1 U411 ( .A(KEYINPUT38), .ZN(n413) );
  XNOR2_X1 U412 ( .A(G101), .B(KEYINPUT71), .ZN(n464) );
  XNOR2_X1 U413 ( .A(n453), .B(n452), .ZN(n465) );
  XNOR2_X1 U414 ( .A(n647), .B(KEYINPUT82), .ZN(n443) );
  AND2_X1 U415 ( .A1(n522), .A2(n423), .ZN(n422) );
  AND2_X1 U416 ( .A1(n664), .A2(n663), .ZN(n469) );
  INV_X1 U417 ( .A(n596), .ZN(n372) );
  NAND2_X1 U418 ( .A1(n411), .A2(n373), .ZN(n410) );
  XNOR2_X1 U419 ( .A(n445), .B(n444), .ZN(n548) );
  INV_X1 U420 ( .A(KEYINPUT8), .ZN(n444) );
  NAND2_X1 U421 ( .A1(n527), .A2(G234), .ZN(n445) );
  AND2_X1 U422 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U423 ( .A1(n620), .A2(n440), .ZN(n436) );
  NOR2_X1 U424 ( .A1(n609), .A2(n608), .ZN(n629) );
  XNOR2_X1 U425 ( .A(n472), .B(n628), .ZN(n471) );
  NOR2_X1 U426 ( .A1(n610), .A2(n515), .ZN(n472) );
  INV_X1 U427 ( .A(KEYINPUT19), .ZN(n455) );
  AND2_X1 U428 ( .A1(n454), .A2(n457), .ZN(n428) );
  NAND2_X1 U429 ( .A1(n515), .A2(KEYINPUT19), .ZN(n457) );
  NAND2_X1 U430 ( .A1(n725), .A2(n724), .ZN(n721) );
  XNOR2_X1 U431 ( .A(G116), .B(G107), .ZN(n493) );
  INV_X1 U432 ( .A(KEYINPUT102), .ZN(n492) );
  XNOR2_X1 U433 ( .A(n506), .B(G134), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n491), .B(n359), .ZN(n416) );
  XNOR2_X1 U435 ( .A(n611), .B(KEYINPUT28), .ZN(n614) );
  XNOR2_X1 U436 ( .A(n636), .B(KEYINPUT111), .ZN(n637) );
  NAND2_X1 U437 ( .A1(n473), .A2(n478), .ZN(n475) );
  XNOR2_X1 U438 ( .A(n531), .B(n500), .ZN(n462) );
  XNOR2_X1 U439 ( .A(KEYINPUT16), .B(G122), .ZN(n500) );
  NOR2_X1 U440 ( .A1(n698), .A2(n358), .ZN(n442) );
  XNOR2_X1 U441 ( .A(n391), .B(n390), .ZN(n616) );
  INV_X1 U442 ( .A(KEYINPUT83), .ZN(n390) );
  OR2_X2 U443 ( .A1(n679), .A2(n569), .ZN(n374) );
  INV_X1 U444 ( .A(KEYINPUT86), .ZN(n441) );
  INV_X1 U445 ( .A(n391), .ZN(n715) );
  INV_X1 U446 ( .A(G237), .ZN(n511) );
  INV_X1 U447 ( .A(n525), .ZN(n401) );
  NAND2_X1 U448 ( .A1(n382), .A2(G902), .ZN(n380) );
  NAND2_X1 U449 ( .A1(n425), .A2(n421), .ZN(n402) );
  AND2_X1 U450 ( .A1(n427), .A2(n524), .ZN(n426) );
  XNOR2_X1 U451 ( .A(G146), .B(G137), .ZN(n539) );
  XNOR2_X1 U452 ( .A(n370), .B(n526), .ZN(n544) );
  XNOR2_X1 U453 ( .A(KEYINPUT4), .B(G131), .ZN(n526) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n516) );
  INV_X1 U455 ( .A(n634), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n383), .B(n354), .ZN(n582) );
  OR2_X1 U457 ( .A1(n667), .A2(G902), .ZN(n383) );
  NOR2_X1 U458 ( .A1(n522), .A2(n423), .ZN(n418) );
  INV_X1 U459 ( .A(n422), .ZN(n420) );
  INV_X1 U460 ( .A(n402), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n558), .B(n560), .ZN(n449) );
  INV_X1 U462 ( .A(KEYINPUT45), .ZN(n406) );
  XNOR2_X1 U463 ( .A(G137), .B(G140), .ZN(n547) );
  XNOR2_X1 U464 ( .A(G119), .B(G110), .ZN(n551) );
  XNOR2_X1 U465 ( .A(G113), .B(G131), .ZN(n487) );
  INV_X1 U466 ( .A(G140), .ZN(n490) );
  XNOR2_X1 U467 ( .A(n353), .B(n488), .ZN(n459) );
  XNOR2_X1 U468 ( .A(n489), .B(n486), .ZN(n460) );
  XOR2_X1 U469 ( .A(G101), .B(G146), .Z(n529) );
  NOR2_X1 U470 ( .A1(n700), .A2(n477), .ZN(n476) );
  INV_X1 U471 ( .A(n700), .ZN(n621) );
  AND2_X1 U472 ( .A1(n471), .A2(n470), .ZN(n630) );
  INV_X1 U473 ( .A(n629), .ZN(n470) );
  XNOR2_X1 U474 ( .A(n447), .B(KEYINPUT80), .ZN(n646) );
  NOR2_X1 U475 ( .A1(n355), .A2(n612), .ZN(n446) );
  XNOR2_X1 U476 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U477 ( .A(KEYINPUT100), .ZN(n581) );
  XNOR2_X1 U478 ( .A(n417), .B(n415), .ZN(n758) );
  XNOR2_X1 U479 ( .A(n495), .B(n494), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n385), .B(n384), .ZN(n667) );
  XNOR2_X1 U481 ( .A(n460), .B(n461), .ZN(n384) );
  XNOR2_X1 U482 ( .A(n766), .B(n459), .ZN(n385) );
  XNOR2_X1 U483 ( .A(n487), .B(n490), .ZN(n461) );
  BUF_X1 U484 ( .A(n752), .Z(n761) );
  XNOR2_X1 U485 ( .A(n601), .B(n510), .ZN(n674) );
  AND2_X1 U486 ( .A1(n670), .A2(G953), .ZN(n765) );
  NAND2_X1 U487 ( .A1(n614), .A2(n613), .ZN(n639) );
  XNOR2_X1 U488 ( .A(n483), .B(n482), .ZN(n781) );
  INV_X1 U489 ( .A(KEYINPUT40), .ZN(n482) );
  NAND2_X1 U490 ( .A1(n474), .A2(n475), .ZN(n483) );
  AND2_X1 U491 ( .A1(n480), .A2(n476), .ZN(n474) );
  INV_X1 U492 ( .A(n724), .ZN(n451) );
  XOR2_X1 U493 ( .A(KEYINPUT99), .B(G122), .Z(n353) );
  INV_X1 U494 ( .A(n725), .ZN(n448) );
  XOR2_X1 U495 ( .A(G475), .B(KEYINPUT13), .Z(n354) );
  XNOR2_X1 U496 ( .A(n375), .B(KEYINPUT35), .ZN(n778) );
  AND2_X1 U497 ( .A1(n428), .A2(n427), .ZN(n355) );
  AND2_X1 U498 ( .A1(n443), .A2(n442), .ZN(n356) );
  OR2_X1 U499 ( .A1(n596), .A2(n595), .ZN(n357) );
  AND2_X1 U500 ( .A1(n715), .A2(KEYINPUT47), .ZN(n358) );
  XOR2_X1 U501 ( .A(G122), .B(KEYINPUT101), .Z(n359) );
  NOR2_X1 U502 ( .A1(n658), .A2(n768), .ZN(n360) );
  AND2_X1 U503 ( .A1(n724), .A2(n525), .ZN(n361) );
  AND2_X1 U504 ( .A1(n480), .A2(n479), .ZN(n362) );
  INV_X1 U505 ( .A(G902), .ZN(n378) );
  AND2_X1 U506 ( .A1(n711), .A2(n455), .ZN(n363) );
  INV_X1 U507 ( .A(KEYINPUT108), .ZN(n440) );
  XOR2_X1 U508 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n364) );
  XNOR2_X1 U509 ( .A(n545), .B(n462), .ZN(n601) );
  NAND2_X1 U510 ( .A1(KEYINPUT84), .A2(n662), .ZN(n365) );
  XNOR2_X2 U511 ( .A(n632), .B(KEYINPUT76), .ZN(n645) );
  NAND2_X1 U512 ( .A1(n614), .A2(n446), .ZN(n447) );
  NAND2_X1 U513 ( .A1(n518), .A2(G902), .ZN(n367) );
  BUF_X2 U514 ( .A(n610), .Z(n368) );
  NAND2_X1 U515 ( .A1(n393), .A2(n403), .ZN(n392) );
  NAND2_X1 U516 ( .A1(n357), .A2(n369), .ZN(n411) );
  NAND2_X1 U517 ( .A1(n596), .A2(n441), .ZN(n369) );
  XNOR2_X1 U518 ( .A(n416), .B(n370), .ZN(n415) );
  NAND2_X1 U519 ( .A1(n371), .A2(KEYINPUT44), .ZN(n409) );
  NAND2_X1 U520 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U521 ( .A(n778), .ZN(n373) );
  XNOR2_X2 U522 ( .A(n374), .B(n570), .ZN(n596) );
  NAND2_X1 U523 ( .A1(n575), .A2(n642), .ZN(n375) );
  NAND2_X1 U524 ( .A1(n754), .A2(n382), .ZN(n381) );
  INV_X1 U525 ( .A(n535), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U527 ( .A(n412), .B(KEYINPUT46), .ZN(n389) );
  NAND2_X1 U528 ( .A1(n403), .A2(n405), .ZN(n573) );
  NAND2_X1 U529 ( .A1(n396), .A2(n392), .ZN(n566) );
  NAND2_X1 U530 ( .A1(n404), .A2(n361), .ZN(n394) );
  INV_X1 U531 ( .A(n405), .ZN(n395) );
  NAND2_X1 U532 ( .A1(n398), .A2(n401), .ZN(n397) );
  NAND2_X1 U533 ( .A1(n399), .A2(n405), .ZN(n398) );
  NOR2_X1 U534 ( .A1(n634), .A2(n451), .ZN(n399) );
  NAND2_X1 U535 ( .A1(n402), .A2(n401), .ZN(n400) );
  NOR2_X2 U536 ( .A1(n419), .A2(n418), .ZN(n405) );
  XNOR2_X2 U537 ( .A(n407), .B(n406), .ZN(n658) );
  INV_X1 U538 ( .A(n428), .ZN(n424) );
  NOR2_X1 U539 ( .A1(n768), .A2(n365), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n638), .B(n637), .ZN(n736) );
  NOR2_X1 U541 ( .A1(n777), .A2(n781), .ZN(n412) );
  XNOR2_X2 U542 ( .A(n654), .B(n413), .ZN(n635) );
  NOR2_X1 U543 ( .A1(n427), .A2(n420), .ZN(n419) );
  NAND2_X1 U544 ( .A1(n424), .A2(n422), .ZN(n421) );
  INV_X1 U545 ( .A(n524), .ZN(n423) );
  NAND2_X1 U546 ( .A1(n426), .A2(n428), .ZN(n425) );
  NAND2_X1 U547 ( .A1(n429), .A2(n662), .ZN(n430) );
  INV_X1 U548 ( .A(n768), .ZN(n429) );
  OR2_X1 U549 ( .A1(n658), .A2(n430), .ZN(n661) );
  NAND2_X1 U550 ( .A1(n432), .A2(n431), .ZN(n664) );
  INV_X1 U551 ( .A(n658), .ZN(n432) );
  NAND2_X1 U552 ( .A1(n627), .A2(n356), .ZN(n433) );
  NAND2_X1 U553 ( .A1(n435), .A2(n434), .ZN(n622) );
  NAND2_X1 U554 ( .A1(n439), .A2(n576), .ZN(n434) );
  XNOR2_X2 U555 ( .A(n368), .B(KEYINPUT6), .ZN(n576) );
  NAND2_X1 U556 ( .A1(n438), .A2(n440), .ZN(n437) );
  NOR2_X1 U557 ( .A1(n620), .A2(n440), .ZN(n439) );
  NAND2_X1 U558 ( .A1(n469), .A2(n468), .ZN(n467) );
  INV_X1 U559 ( .A(n633), .ZN(n456) );
  NAND2_X1 U560 ( .A1(n633), .A2(KEYINPUT19), .ZN(n454) );
  NAND2_X1 U561 ( .A1(n643), .A2(n711), .ZN(n623) );
  NOR2_X1 U562 ( .A1(n758), .A2(G902), .ZN(n458) );
  XNOR2_X2 U563 ( .A(G110), .B(G107), .ZN(n463) );
  XNOR2_X2 U564 ( .A(n513), .B(n512), .ZN(n633) );
  NAND2_X1 U565 ( .A1(n466), .A2(n665), .ZN(n681) );
  XNOR2_X1 U566 ( .A(n467), .B(KEYINPUT64), .ZN(n466) );
  NAND2_X1 U567 ( .A1(n661), .A2(n660), .ZN(n468) );
  INV_X1 U568 ( .A(n368), .ZN(n728) );
  INV_X1 U569 ( .A(n645), .ZN(n473) );
  NAND2_X1 U570 ( .A1(n645), .A2(n481), .ZN(n480) );
  NAND2_X1 U571 ( .A1(n362), .A2(n475), .ZN(n655) );
  INV_X1 U572 ( .A(n479), .ZN(n477) );
  NOR2_X1 U573 ( .A1(n635), .A2(n481), .ZN(n478) );
  NAND2_X1 U574 ( .A1(n635), .A2(n481), .ZN(n479) );
  INV_X1 U575 ( .A(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U576 ( .A(n484), .B(n544), .ZN(n683) );
  XNOR2_X1 U577 ( .A(n543), .B(n545), .ZN(n484) );
  XNOR2_X1 U578 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X2 U579 ( .A(n568), .B(n567), .ZN(n679) );
  XNOR2_X2 U580 ( .A(n504), .B(KEYINPUT10), .ZN(n766) );
  XOR2_X2 U581 ( .A(G146), .B(G125), .Z(n504) );
  XOR2_X1 U582 ( .A(n653), .B(KEYINPUT109), .Z(n485) );
  INV_X1 U583 ( .A(KEYINPUT84), .ZN(n660) );
  XNOR2_X1 U584 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U585 ( .A(n557), .B(KEYINPUT93), .ZN(n558) );
  XNOR2_X1 U586 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U587 ( .A(KEYINPUT41), .ZN(n636) );
  XNOR2_X1 U588 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n767), .B(n532), .ZN(n754) );
  XNOR2_X1 U590 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U591 ( .A(G143), .B(G104), .ZN(n486) );
  XOR2_X1 U592 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n489) );
  NOR2_X2 U593 ( .A1(G953), .A2(G237), .ZN(n536) );
  NAND2_X1 U594 ( .A1(G214), .A2(n536), .ZN(n488) );
  XNOR2_X2 U595 ( .A(G143), .B(G128), .ZN(n506) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n491) );
  NAND2_X1 U597 ( .A1(G217), .A2(n548), .ZN(n495) );
  XNOR2_X1 U598 ( .A(KEYINPUT103), .B(G478), .ZN(n496) );
  NAND2_X1 U599 ( .A1(n659), .A2(G234), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n497), .B(KEYINPUT20), .ZN(n556) );
  AND2_X1 U601 ( .A1(n556), .A2(G221), .ZN(n499) );
  XNOR2_X1 U602 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n498) );
  XNOR2_X1 U603 ( .A(n499), .B(n498), .ZN(n724) );
  XNOR2_X1 U604 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n527), .A2(G224), .ZN(n501) );
  XNOR2_X1 U606 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n509) );
  XNOR2_X1 U608 ( .A(KEYINPUT4), .B(KEYINPUT77), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n352), .B(n505), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U611 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U612 ( .A1(n674), .A2(n659), .ZN(n513) );
  NAND2_X1 U613 ( .A1(n378), .A2(n511), .ZN(n514) );
  NAND2_X1 U614 ( .A1(n514), .A2(G210), .ZN(n512) );
  NAND2_X1 U615 ( .A1(n514), .A2(G214), .ZN(n711) );
  INV_X1 U616 ( .A(n711), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(KEYINPUT14), .ZN(n518) );
  NAND2_X1 U618 ( .A1(n518), .A2(G952), .ZN(n517) );
  XOR2_X1 U619 ( .A(KEYINPUT91), .B(n517), .Z(n743) );
  NOR2_X1 U620 ( .A1(n743), .A2(G953), .ZN(n609) );
  INV_X1 U621 ( .A(n609), .ZN(n521) );
  NAND2_X1 U622 ( .A1(G953), .A2(n519), .ZN(n606) );
  OR2_X1 U623 ( .A1(n606), .A2(G898), .ZN(n520) );
  NAND2_X1 U624 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U625 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n523) );
  XNOR2_X1 U626 ( .A(n523), .B(KEYINPUT66), .ZN(n524) );
  XNOR2_X1 U627 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n544), .B(n547), .ZN(n767) );
  NAND2_X1 U629 ( .A1(G227), .A2(n527), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U632 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n534) );
  INV_X1 U633 ( .A(G469), .ZN(n533) );
  AND2_X1 U634 ( .A1(n566), .A2(n722), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n538) );
  NAND2_X1 U636 ( .A1(n536), .A2(G210), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n538), .B(n537), .ZN(n542) );
  XOR2_X1 U638 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n540) );
  XNOR2_X1 U639 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U640 ( .A1(n683), .A2(n378), .ZN(n546) );
  INV_X1 U641 ( .A(G472), .ZN(n680) );
  XNOR2_X1 U642 ( .A(n547), .B(G128), .ZN(n550) );
  NAND2_X1 U643 ( .A1(G221), .A2(n548), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n550), .B(n549), .ZN(n555) );
  XOR2_X1 U645 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n552) );
  XNOR2_X1 U646 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n766), .B(n553), .ZN(n554) );
  XNOR2_X1 U648 ( .A(n554), .B(n555), .ZN(n762) );
  NOR2_X1 U649 ( .A1(n762), .A2(G902), .ZN(n559) );
  NAND2_X1 U650 ( .A1(G217), .A2(n556), .ZN(n557) );
  INV_X1 U651 ( .A(KEYINPUT25), .ZN(n560) );
  AND2_X1 U652 ( .A1(n368), .A2(n448), .ZN(n561) );
  AND2_X1 U653 ( .A1(n577), .A2(n561), .ZN(n569) );
  XOR2_X1 U654 ( .A(G110), .B(n569), .Z(G12) );
  OR2_X1 U655 ( .A1(n722), .A2(n725), .ZN(n564) );
  INV_X1 U656 ( .A(KEYINPUT79), .ZN(n562) );
  XNOR2_X1 U657 ( .A(n576), .B(n562), .ZN(n563) );
  NOR2_X1 U658 ( .A1(n564), .A2(n563), .ZN(n565) );
  AND2_X2 U659 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U660 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n567) );
  INV_X1 U661 ( .A(KEYINPUT87), .ZN(n570) );
  INV_X1 U662 ( .A(KEYINPUT33), .ZN(n572) );
  NAND2_X1 U663 ( .A1(n585), .A2(n576), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n572), .B(n571), .ZN(n718) );
  NOR2_X1 U665 ( .A1(n718), .A2(n573), .ZN(n574) );
  XNOR2_X1 U666 ( .A(n574), .B(KEYINPUT34), .ZN(n575) );
  AND2_X1 U667 ( .A1(n584), .A2(n582), .ZN(n642) );
  AND2_X1 U668 ( .A1(n577), .A2(n438), .ZN(n578) );
  XNOR2_X1 U669 ( .A(n578), .B(KEYINPUT85), .ZN(n579) );
  NOR2_X1 U670 ( .A1(n579), .A2(n448), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n580), .B(KEYINPUT106), .ZN(n782) );
  NAND2_X1 U672 ( .A1(n584), .A2(n583), .ZN(n702) );
  NAND2_X1 U673 ( .A1(n728), .A2(n585), .ZN(n731) );
  NOR2_X1 U674 ( .A1(n573), .A2(n731), .ZN(n587) );
  XNOR2_X1 U675 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n586) );
  XNOR2_X1 U676 ( .A(n587), .B(n586), .ZN(n703) );
  NOR2_X1 U677 ( .A1(n612), .A2(n721), .ZN(n631) );
  NAND2_X1 U678 ( .A1(n631), .A2(n368), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n588), .A2(n573), .ZN(n589) );
  XNOR2_X1 U680 ( .A(KEYINPUT97), .B(n589), .ZN(n690) );
  NAND2_X1 U681 ( .A1(n703), .A2(n690), .ZN(n590) );
  NAND2_X1 U682 ( .A1(n616), .A2(n590), .ZN(n591) );
  XOR2_X1 U683 ( .A(KEYINPUT104), .B(n591), .Z(n592) );
  NOR2_X1 U684 ( .A1(n782), .A2(n592), .ZN(n593) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n594), .A2(KEYINPUT86), .ZN(n595) );
  NOR2_X1 U687 ( .A1(n658), .A2(G953), .ZN(n600) );
  INV_X1 U688 ( .A(G898), .ZN(n602) );
  NAND2_X1 U689 ( .A1(G953), .A2(G224), .ZN(n597) );
  XOR2_X1 U690 ( .A(KEYINPUT61), .B(n597), .Z(n598) );
  NOR2_X1 U691 ( .A1(n602), .A2(n598), .ZN(n599) );
  NOR2_X1 U692 ( .A1(n600), .A2(n599), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n602), .A2(G953), .ZN(n603) );
  NAND2_X1 U694 ( .A1(n601), .A2(n603), .ZN(n604) );
  XNOR2_X1 U695 ( .A(n605), .B(n604), .ZN(G69) );
  NOR2_X1 U696 ( .A1(G900), .A2(n606), .ZN(n607) );
  XOR2_X1 U697 ( .A(KEYINPUT107), .B(n607), .Z(n608) );
  NOR2_X1 U698 ( .A1(n610), .A2(n620), .ZN(n611) );
  INV_X1 U699 ( .A(n612), .ZN(n613) );
  XNOR2_X1 U700 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U702 ( .A(n617), .B(KEYINPUT74), .ZN(n618) );
  XNOR2_X1 U703 ( .A(n619), .B(KEYINPUT73), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n648) );
  NOR2_X1 U705 ( .A1(n648), .A2(n623), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n624), .B(KEYINPUT36), .ZN(n625) );
  INV_X1 U707 ( .A(n722), .ZN(n651) );
  NAND2_X1 U708 ( .A1(n625), .A2(n651), .ZN(n626) );
  XNOR2_X1 U709 ( .A(n626), .B(KEYINPUT113), .ZN(n779) );
  XNOR2_X1 U710 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U712 ( .A(n635), .ZN(n712) );
  NAND2_X1 U713 ( .A1(n712), .A2(n711), .ZN(n714) );
  NOR2_X1 U714 ( .A1(n634), .A2(n714), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n736), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n777) );
  INV_X1 U718 ( .A(n654), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n698) );
  NAND2_X1 U721 ( .A1(n646), .A2(KEYINPUT47), .ZN(n647) );
  INV_X1 U722 ( .A(n648), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n649), .A2(n711), .ZN(n650) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U725 ( .A(KEYINPUT43), .B(n652), .Z(n653) );
  NAND2_X1 U726 ( .A1(n485), .A2(n654), .ZN(n707) );
  NOR2_X1 U727 ( .A1(n702), .A2(n655), .ZN(n705) );
  INV_X1 U728 ( .A(n705), .ZN(n656) );
  AND2_X1 U729 ( .A1(n707), .A2(n656), .ZN(n657) );
  INV_X1 U730 ( .A(n659), .ZN(n662) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n709) );
  OR2_X1 U732 ( .A1(n659), .A2(n709), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n360), .A2(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n752), .A2(G475), .ZN(n669) );
  XNOR2_X1 U735 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n669), .B(n668), .ZN(n671) );
  INV_X1 U737 ( .A(G952), .ZN(n670) );
  NOR2_X2 U738 ( .A1(n671), .A2(n765), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U740 ( .A1(n752), .A2(G210), .ZN(n676) );
  XNOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X2 U744 ( .A1(n677), .A2(n765), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U746 ( .A(n679), .B(G119), .Z(G21) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n685) );
  XNOR2_X1 U748 ( .A(KEYINPUT90), .B(KEYINPUT62), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n686), .A2(n765), .ZN(n688) );
  XOR2_X1 U752 ( .A(KEYINPUT114), .B(KEYINPUT63), .Z(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(G57) );
  NOR2_X1 U754 ( .A1(n700), .A2(n690), .ZN(n689) );
  XOR2_X1 U755 ( .A(G104), .B(n689), .Z(G6) );
  NOR2_X1 U756 ( .A1(n690), .A2(n702), .ZN(n694) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n692) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U759 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n694), .B(n693), .ZN(G9) );
  NOR2_X1 U761 ( .A1(n646), .A2(n702), .ZN(n696) );
  XNOR2_X1 U762 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(G128), .B(n697), .ZN(G30) );
  XOR2_X1 U765 ( .A(G143), .B(n698), .Z(G45) );
  NOR2_X1 U766 ( .A1(n646), .A2(n700), .ZN(n699) );
  XOR2_X1 U767 ( .A(G146), .B(n699), .Z(G48) );
  NOR2_X1 U768 ( .A1(n703), .A2(n700), .ZN(n701) );
  XOR2_X1 U769 ( .A(G113), .B(n701), .Z(G15) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U771 ( .A(G116), .B(n704), .Z(G18) );
  XNOR2_X1 U772 ( .A(G134), .B(n705), .ZN(n706) );
  XNOR2_X1 U773 ( .A(n706), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U774 ( .A(n707), .B(G140), .ZN(n708) );
  XNOR2_X1 U775 ( .A(KEYINPUT118), .B(n708), .ZN(G42) );
  NOR2_X1 U776 ( .A1(n360), .A2(KEYINPUT81), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(n709), .ZN(n748) );
  NOR2_X1 U778 ( .A1(n736), .A2(n718), .ZN(n746) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U780 ( .A1(n634), .A2(n713), .ZN(n717) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n719) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n739) );
  XNOR2_X1 U784 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n720) );
  XNOR2_X1 U785 ( .A(n720), .B(KEYINPUT51), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U787 ( .A(n723), .B(KEYINPUT50), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U789 ( .A(KEYINPUT49), .B(n726), .Z(n727) );
  NOR2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U791 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U793 ( .A(n734), .B(n733), .Z(n735) );
  NOR2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U795 ( .A(KEYINPUT121), .B(n737), .Z(n738) );
  NOR2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n742) );
  XOR2_X1 U797 ( .A(KEYINPUT52), .B(KEYINPUT123), .Z(n740) );
  XNOR2_X1 U798 ( .A(KEYINPUT122), .B(n740), .ZN(n741) );
  XNOR2_X1 U799 ( .A(n742), .B(n741), .ZN(n744) );
  NOR2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U801 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U803 ( .A(KEYINPUT124), .B(n749), .ZN(n750) );
  NOR2_X1 U804 ( .A1(n750), .A2(G953), .ZN(n751) );
  XNOR2_X1 U805 ( .A(n751), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U806 ( .A1(n761), .A2(G469), .ZN(n756) );
  XOR2_X1 U807 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n753) );
  NOR2_X1 U808 ( .A1(n765), .A2(n757), .ZN(G54) );
  NAND2_X1 U809 ( .A1(n761), .A2(G478), .ZN(n759) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n765), .A2(n760), .ZN(G63) );
  NAND2_X1 U812 ( .A1(n761), .A2(G217), .ZN(n763) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U814 ( .A1(n765), .A2(n764), .ZN(G66) );
  XNOR2_X1 U815 ( .A(n767), .B(n766), .ZN(n770) );
  XOR2_X1 U816 ( .A(n770), .B(n768), .Z(n769) );
  NOR2_X1 U817 ( .A1(G953), .A2(n769), .ZN(n775) );
  XNOR2_X1 U818 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(G953), .ZN(n773) );
  XOR2_X1 U821 ( .A(KEYINPUT126), .B(n773), .Z(n774) );
  NOR2_X1 U822 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U823 ( .A(KEYINPUT127), .B(n776), .ZN(G72) );
  XOR2_X1 U824 ( .A(G137), .B(n777), .Z(G39) );
  XOR2_X1 U825 ( .A(G122), .B(n778), .Z(G24) );
  XNOR2_X1 U826 ( .A(G125), .B(n779), .ZN(n780) );
  XNOR2_X1 U827 ( .A(n780), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U828 ( .A(n781), .B(G131), .Z(G33) );
  XOR2_X1 U829 ( .A(G101), .B(n782), .Z(G3) );
endmodule

