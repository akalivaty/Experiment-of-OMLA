

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  OR2_X1 U324 ( .A1(n394), .A2(n393), .ZN(n395) );
  NOR2_X1 U325 ( .A1(n531), .A2(n451), .ZN(n452) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n292) );
  XOR2_X1 U327 ( .A(n364), .B(n363), .Z(n293) );
  XOR2_X1 U328 ( .A(KEYINPUT105), .B(n396), .Z(n294) );
  INV_X1 U329 ( .A(n578), .ZN(n389) );
  XNOR2_X1 U330 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n328), .B(n327), .ZN(n333) );
  XNOR2_X1 U332 ( .A(n365), .B(n293), .ZN(n366) );
  XNOR2_X1 U333 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U334 ( .A(KEYINPUT118), .B(n452), .ZN(n569) );
  XOR2_X1 U335 ( .A(KEYINPUT41), .B(n583), .Z(n555) );
  XNOR2_X1 U336 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XNOR2_X1 U338 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n295), .B(G183GAT), .ZN(n296) );
  XOR2_X1 U340 ( .A(n296), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n410) );
  XOR2_X1 U343 ( .A(G134GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U350 ( .A(G15GAT), .B(KEYINPUT64), .Z(n306) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(n307), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n410), .B(n310), .ZN(n314) );
  XOR2_X1 U356 ( .A(KEYINPUT82), .B(G127GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(G113GAT), .B(n313), .Z(n429) );
  XOR2_X1 U360 ( .A(n314), .B(n429), .Z(n531) );
  XOR2_X1 U361 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n316) );
  XNOR2_X1 U362 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n315) );
  XOR2_X1 U363 ( .A(n316), .B(n315), .Z(n335) );
  INV_X1 U364 ( .A(KEYINPUT69), .ZN(n317) );
  NAND2_X1 U365 ( .A1(n317), .A2(G57GAT), .ZN(n320) );
  INV_X1 U366 ( .A(G57GAT), .ZN(n318) );
  NAND2_X1 U367 ( .A1(n318), .A2(KEYINPUT69), .ZN(n319) );
  NAND2_X1 U368 ( .A1(n320), .A2(n319), .ZN(n322) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n351) );
  XOR2_X1 U371 ( .A(G99GAT), .B(G85GAT), .Z(n357) );
  XNOR2_X1 U372 ( .A(n351), .B(n357), .ZN(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n324) );
  XNOR2_X1 U374 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n326) );
  AND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n329), .B(G148GAT), .ZN(n435) );
  XOR2_X1 U379 ( .A(G64GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n405) );
  XOR2_X1 U382 ( .A(n435), .B(n405), .Z(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n478) );
  INV_X1 U385 ( .A(n478), .ZN(n583) );
  XOR2_X1 U386 ( .A(G64GAT), .B(G127GAT), .Z(n337) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n473) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XOR2_X1 U390 ( .A(n436), .B(G78GAT), .Z(n339) );
  XOR2_X1 U391 ( .A(G15GAT), .B(G1GAT), .Z(n384) );
  XNOR2_X1 U392 ( .A(n384), .B(G211GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n341) );
  XNOR2_X1 U395 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n340) );
  XOR2_X1 U396 ( .A(n341), .B(n340), .Z(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n345) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n347) );
  INV_X1 U400 ( .A(KEYINPUT78), .ZN(n346) );
  NAND2_X1 U401 ( .A1(n347), .A2(n346), .ZN(n350) );
  INV_X1 U402 ( .A(n347), .ZN(n348) );
  NAND2_X1 U403 ( .A1(n348), .A2(KEYINPUT78), .ZN(n349) );
  NAND2_X1 U404 ( .A1(n350), .A2(n349), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n351), .B(KEYINPUT14), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n472) );
  XNOR2_X1 U407 ( .A(n473), .B(n472), .ZN(n491) );
  XOR2_X1 U408 ( .A(G29GAT), .B(G43GAT), .Z(n355) );
  XNOR2_X1 U409 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n386) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n356), .B(G162GAT), .ZN(n439) );
  XNOR2_X1 U413 ( .A(n386), .B(n439), .ZN(n369) );
  XOR2_X1 U414 ( .A(G134GAT), .B(KEYINPUT77), .Z(n415) );
  XOR2_X1 U415 ( .A(n357), .B(n415), .Z(n359) );
  NAND2_X1 U416 ( .A1(G232GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n367) );
  XOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .Z(n403) );
  XOR2_X1 U419 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n361) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n403), .B(n362), .ZN(n365) );
  XOR2_X1 U423 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n364) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(G92GAT), .ZN(n363) );
  XOR2_X1 U425 ( .A(n369), .B(n368), .Z(n568) );
  XOR2_X1 U426 ( .A(n568), .B(KEYINPUT36), .Z(n589) );
  NOR2_X1 U427 ( .A1(n491), .A2(n589), .ZN(n370) );
  XOR2_X1 U428 ( .A(KEYINPUT45), .B(n370), .Z(n371) );
  NOR2_X1 U429 ( .A1(n583), .A2(n371), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n372), .B(KEYINPUT106), .ZN(n390) );
  XOR2_X1 U431 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n374) );
  NAND2_X1 U432 ( .A1(G229GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U434 ( .A(n375), .B(KEYINPUT66), .Z(n383) );
  XOR2_X1 U435 ( .A(G141GAT), .B(G197GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(G36GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U438 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n379) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G113GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U443 ( .A(n385), .B(n384), .Z(n388) );
  XOR2_X1 U444 ( .A(G169GAT), .B(G8GAT), .Z(n406) );
  XNOR2_X1 U445 ( .A(n386), .B(n406), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n578) );
  AND2_X1 U447 ( .A1(n390), .A2(n389), .ZN(n397) );
  NAND2_X1 U448 ( .A1(n578), .A2(n555), .ZN(n392) );
  XOR2_X1 U449 ( .A(KEYINPUT104), .B(KEYINPUT46), .Z(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n394) );
  INV_X1 U451 ( .A(n568), .ZN(n474) );
  NAND2_X1 U452 ( .A1(n491), .A2(n474), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n395), .B(KEYINPUT47), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n397), .A2(n294), .ZN(n398) );
  XOR2_X1 U455 ( .A(KEYINPUT48), .B(n398), .Z(n530) );
  XOR2_X1 U456 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n445) );
  XOR2_X1 U459 ( .A(KEYINPUT92), .B(n445), .Z(n402) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U462 ( .A(n404), .B(n403), .Z(n408) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U465 ( .A(n410), .B(n409), .Z(n522) );
  INV_X1 U466 ( .A(n522), .ZN(n459) );
  AND2_X1 U467 ( .A1(n530), .A2(n459), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n411), .B(n292), .ZN(n432) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G162GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U475 ( .A(n418), .B(KEYINPUT1), .Z(n421) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n419), .B(KEYINPUT2), .ZN(n444) );
  XNOR2_X1 U478 ( .A(n444), .B(KEYINPUT91), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT6), .B(G57GAT), .Z(n423) );
  XNOR2_X1 U481 ( .A(G1GAT), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n520) );
  INV_X1 U489 ( .A(n520), .ZN(n469) );
  NOR2_X1 U490 ( .A1(n432), .A2(n469), .ZN(n575) );
  XOR2_X1 U491 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n434) );
  XNOR2_X1 U492 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U494 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U495 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n443) );
  XOR2_X1 U497 ( .A(n439), .B(KEYINPUT24), .Z(n441) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U500 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n463) );
  NAND2_X1 U504 ( .A1(n575), .A2(n463), .ZN(n450) );
  XOR2_X1 U505 ( .A(n450), .B(KEYINPUT55), .Z(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT99), .B(n555), .ZN(n507) );
  INV_X1 U507 ( .A(n507), .ZN(n537) );
  NAND2_X1 U508 ( .A1(n569), .A2(n537), .ZN(n456) );
  XOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n453) );
  INV_X1 U511 ( .A(n531), .ZN(n462) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n522), .ZN(n465) );
  NOR2_X1 U513 ( .A1(n520), .A2(n465), .ZN(n529) );
  XNOR2_X1 U514 ( .A(n463), .B(KEYINPUT28), .ZN(n528) );
  NAND2_X1 U515 ( .A1(n529), .A2(n528), .ZN(n457) );
  XOR2_X1 U516 ( .A(KEYINPUT93), .B(n457), .Z(n458) );
  NOR2_X1 U517 ( .A1(n462), .A2(n458), .ZN(n471) );
  NAND2_X1 U518 ( .A1(n462), .A2(n459), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n463), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT25), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U522 ( .A(n464), .B(KEYINPUT26), .Z(n574) );
  NOR2_X1 U523 ( .A1(n465), .A2(n574), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n489) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n476) );
  XOR2_X1 U528 ( .A(n473), .B(n472), .Z(n586) );
  NAND2_X1 U529 ( .A1(n586), .A2(n474), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U531 ( .A1(n489), .A2(n477), .ZN(n508) );
  NAND2_X1 U532 ( .A1(n478), .A2(n578), .ZN(n479) );
  XOR2_X1 U533 ( .A(KEYINPUT74), .B(n479), .Z(n493) );
  NAND2_X1 U534 ( .A1(n508), .A2(n493), .ZN(n487) );
  NOR2_X1 U535 ( .A1(n520), .A2(n487), .ZN(n481) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U538 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U539 ( .A1(n522), .A2(n487), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U542 ( .A1(n531), .A2(n487), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U545 ( .A1(n528), .A2(n487), .ZN(n488) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  NOR2_X1 U547 ( .A1(n489), .A2(n589), .ZN(n490) );
  NAND2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(KEYINPUT37), .ZN(n519) );
  NAND2_X1 U550 ( .A1(n493), .A2(n519), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(KEYINPUT38), .ZN(n503) );
  NOR2_X1 U552 ( .A1(n503), .A2(n520), .ZN(n498) );
  XOR2_X1 U553 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n496) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n522), .A2(n503), .ZN(n499) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U559 ( .A1(n503), .A2(n531), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT98), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n502), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n528), .ZN(n504) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT100), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n510) );
  NOR2_X1 U568 ( .A1(n578), .A2(n507), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n518), .A2(n508), .ZN(n513) );
  NOR2_X1 U570 ( .A1(n520), .A2(n513), .ZN(n509) );
  XOR2_X1 U571 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n522), .A2(n513), .ZN(n511) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n531), .A2(n513), .ZN(n512) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n528), .ZN(n517) );
  XOR2_X1 U577 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n515) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT102), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n518), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n520), .A2(n525), .ZN(n521) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n522), .A2(n525), .ZN(n523) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n525), .ZN(n524) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n528), .A2(n525), .ZN(n526) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT108), .ZN(n536) );
  INV_X1 U592 ( .A(n528), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n548) );
  NOR2_X1 U594 ( .A1(n531), .A2(n548), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT107), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n578), .A2(n545), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT110), .Z(n539) );
  NAND2_X1 U600 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT109), .Z(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT111), .Z(n543) );
  NAND2_X1 U605 ( .A1(n545), .A2(n586), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U609 ( .A1(n545), .A2(n568), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT113), .Z(n551) );
  NOR2_X1 U612 ( .A1(n548), .A2(n574), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT112), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n578), .A2(n559), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n553) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT52), .B(n554), .Z(n557) );
  NAND2_X1 U620 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n586), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n568), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(KEYINPUT116), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  XOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U628 ( .A1(n578), .A2(n569), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U631 ( .A1(n586), .A2(n569), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(n567), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n582) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .Z(n580) );
  INV_X1 U642 ( .A(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(KEYINPUT124), .B(n577), .ZN(n590) );
  INV_X1 U645 ( .A(n590), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n578), .A2(n587), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U648 ( .A(n582), .B(n581), .Z(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U650 ( .A1(n587), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

