//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G475), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT18), .A2(G131), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(KEYINPUT91), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT91), .B(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n190), .B1(new_n197), .B2(KEYINPUT92), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(new_n193), .ZN(new_n199));
  NOR2_X1   g013(.A1(G237), .A2(G953), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n200), .A2(G214), .B1(new_n201), .B2(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT93), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(new_n204), .B2(KEYINPUT92), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n203), .A2(KEYINPUT93), .A3(new_n190), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n206), .A3(G125), .ZN(new_n218));
  OAI211_X1 g032(.A(G146), .B(new_n218), .C1(new_n210), .C2(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n210), .B2(new_n217), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n212), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT95), .B1(new_n203), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n197), .A2(new_n224), .A3(G131), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n219), .B(new_n221), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n203), .A2(KEYINPUT94), .A3(new_n222), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n197), .B2(G131), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n223), .A2(new_n229), .A3(new_n225), .A4(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT17), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n216), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G113), .B(G122), .ZN(new_n235));
  INV_X1    g049(.A(G104), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(new_n216), .C1(new_n228), .C2(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n189), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n219), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n210), .B(KEYINPUT19), .Z(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n212), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n232), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT96), .A3(new_n216), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n238), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT96), .B1(new_n247), .B2(new_n216), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n240), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G475), .A2(G902), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n216), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n238), .A3(new_n248), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT97), .B1(new_n257), .B2(new_n240), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(new_n258), .B2(KEYINPUT20), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n251), .A2(KEYINPUT97), .A3(new_n260), .A4(new_n252), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n243), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(G234), .A2(G237), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n263), .A2(G952), .A3(new_n192), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n263), .A2(G902), .A3(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT21), .B(G898), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(G116), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT14), .A3(G122), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(G122), .ZN(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(G122), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(G107), .B(new_n270), .C1(new_n274), .C2(KEYINPUT14), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n194), .A2(G128), .ZN(new_n278));
  OR2_X1    g092(.A1(KEYINPUT66), .A2(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT66), .A2(G128), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n281), .B2(new_n194), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n275), .A2(new_n277), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G217), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n187), .A2(new_n287), .A3(G953), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n281), .A2(new_n194), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT98), .B(KEYINPUT13), .Z(new_n290));
  OAI21_X1  g104(.A(G134), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(new_n282), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n282), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n274), .B(new_n276), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n286), .B(new_n288), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n288), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n293), .B2(new_n292), .ZN(new_n298));
  INV_X1    g112(.A(new_n286), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT99), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT99), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n242), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT100), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n304), .B(new_n310), .Z(new_n311));
  NAND3_X1  g125(.A1(new_n262), .A2(new_n268), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT101), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n262), .A2(KEYINPUT101), .A3(new_n268), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT11), .B1(new_n283), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n317), .A3(G134), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(new_n222), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n212), .A2(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n194), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n327), .A2(KEYINPUT84), .ZN(new_n328));
  OAI21_X1  g142(.A(G128), .B1(new_n327), .B2(KEYINPUT84), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G128), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(KEYINPUT1), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n324), .A3(new_n325), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT65), .ZN(new_n334));
  XNOR2_X1  g148(.A(G143), .B(G146), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n276), .A2(G104), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n236), .A2(G107), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n236), .B2(G107), .ZN(new_n344));
  AOI21_X1  g158(.A(G101), .B1(new_n236), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n276), .A3(G104), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(KEYINPUT83), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n343), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(KEYINPUT66), .A2(G128), .ZN(new_n355));
  NOR2_X1   g169(.A1(KEYINPUT66), .A2(G128), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G143), .B2(new_n212), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n326), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n336), .B1(new_n335), .B2(new_n332), .ZN(new_n361));
  AND4_X1   g175(.A1(new_n336), .A2(new_n332), .A3(new_n324), .A4(new_n325), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n352), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT12), .B(new_n323), .C1(new_n354), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT85), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n353), .B1(new_n363), .B2(new_n352), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT12), .A4(new_n323), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n323), .B1(new_n354), .B2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n353), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n344), .A2(new_n347), .A3(new_n342), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n376), .A2(new_n377), .A3(G101), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n350), .A2(new_n351), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n376), .B2(G101), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n335), .A2(KEYINPUT0), .A3(G128), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G128), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n335), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n322), .B(G131), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n352), .A2(new_n363), .A3(KEYINPUT10), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n375), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n373), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G110), .B(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n192), .A2(G227), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n375), .A2(new_n386), .A3(new_n388), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n323), .ZN(new_n395));
  INV_X1    g209(.A(new_n393), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n390), .A2(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G469), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n373), .A2(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n393), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G469), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n242), .ZN(new_n405));
  NAND2_X1  g219(.A1(G469), .A2(G902), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n411), .A3(G119), .ZN(new_n412));
  INV_X1    g226(.A(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G116), .ZN(new_n414));
  INV_X1    g228(.A(G113), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT2), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G113), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n412), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n412), .B2(new_n414), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n408), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(new_n414), .ZN(new_n423));
  INV_X1    g237(.A(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n414), .A3(new_n419), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(KEYINPUT68), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n381), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n412), .A2(KEYINPUT5), .A3(new_n414), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n415), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n420), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n352), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n428), .A2(new_n381), .B1(new_n352), .B2(new_n433), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n437), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT86), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n384), .A2(G125), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(G125), .B2(new_n363), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT87), .B(G224), .Z(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n446), .B(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n437), .B1(new_n441), .B2(new_n438), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n435), .A2(new_n439), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT88), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n444), .A2(new_n452), .A3(new_n455), .A4(new_n449), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(new_n447), .B2(G953), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n446), .B(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n441), .B2(new_n438), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n438), .B(KEYINPUT8), .Z(new_n460));
  INV_X1    g274(.A(new_n352), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n433), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n432), .B(KEYINPUT90), .Z(new_n463));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n430), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n430), .A2(new_n464), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(new_n426), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n459), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n456), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G210), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n454), .A2(new_n472), .A3(new_n456), .A4(new_n470), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G214), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AND4_X1   g293(.A1(new_n188), .A2(new_n316), .A3(new_n407), .A4(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT23), .A2(G119), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT23), .A2(G119), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(G128), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n357), .B2(new_n486), .ZN(new_n487));
  NOR4_X1   g301(.A1(new_n355), .A2(new_n356), .A3(new_n482), .A4(KEYINPUT78), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G110), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n221), .A2(new_n219), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n413), .B1(new_n279), .B2(new_n280), .ZN(new_n492));
  NOR2_X1   g306(.A1(G119), .A2(G128), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT77), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT77), .ZN(new_n495));
  INV_X1    g309(.A(new_n493), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n496), .C1(new_n357), .C2(new_n413), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G110), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n490), .B(new_n491), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n499), .A3(new_n497), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(new_n484), .C1(new_n487), .C2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n219), .A2(new_n213), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT79), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n508), .B(new_n505), .C1(new_n501), .C2(new_n503), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n500), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT80), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n500), .B(new_n514), .C1(new_n507), .C2(new_n509), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n242), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(KEYINPUT25), .A3(new_n242), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n287), .B1(G234), .B2(new_n242), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n481), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT81), .B(new_n525), .C1(new_n520), .C2(new_n521), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n516), .A2(new_n517), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n523), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n200), .A2(G210), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT27), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT26), .B(G101), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT64), .B1(new_n317), .B2(G134), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT64), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n283), .A3(G137), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n317), .A2(G134), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G131), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n319), .A2(new_n321), .ZN(new_n545));
  INV_X1    g359(.A(new_n318), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n222), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n323), .A2(new_n385), .B1(new_n548), .B2(new_n363), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n422), .A2(new_n427), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT28), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT72), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT69), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n281), .A2(new_n327), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n334), .A2(new_n337), .B1(new_n554), .B2(new_n326), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n544), .A2(new_n547), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n387), .A2(new_n384), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n557), .B2(new_n428), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT69), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n560), .A3(new_n428), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n552), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n563));
  AOI211_X1 g377(.A(new_n538), .B(new_n551), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n323), .A2(new_n385), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n548), .A2(new_n363), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n550), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n538), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n533), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n558), .A2(new_n559), .ZN(new_n576));
  INV_X1    g390(.A(new_n570), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n569), .B1(new_n567), .B2(new_n568), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n428), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT29), .B1(new_n580), .B2(new_n538), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n562), .A2(new_n563), .ZN(new_n582));
  INV_X1    g396(.A(new_n551), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n537), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT73), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n558), .B(new_n559), .C1(new_n550), .C2(new_n549), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n551), .B1(new_n586), .B2(KEYINPUT28), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n538), .A2(new_n573), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n575), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n590), .A2(KEYINPUT74), .A3(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT74), .B1(new_n590), .B2(G472), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n563), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n557), .A2(new_n560), .A3(new_n428), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n560), .B1(new_n557), .B2(new_n428), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n594), .B1(new_n576), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n538), .B1(new_n598), .B2(new_n551), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n558), .A2(new_n559), .A3(new_n537), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(KEYINPUT70), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n558), .A2(new_n559), .A3(new_n602), .A4(new_n537), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n579), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT31), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(KEYINPUT70), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT31), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n579), .A4(new_n603), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n599), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(G472), .A3(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT75), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n551), .B1(new_n562), .B2(new_n563), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n608), .B1(new_n537), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n603), .A2(new_n579), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n607), .B1(new_n618), .B2(new_n606), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n615), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n610), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n609), .A2(KEYINPUT75), .A3(new_n611), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n614), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT76), .B1(new_n593), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n590), .A2(G472), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT74), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n590), .A2(KEYINPUT74), .A3(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n614), .A2(new_n622), .A3(new_n621), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT76), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n532), .B1(new_n624), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT82), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT82), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n635), .B(new_n532), .C1(new_n624), .C2(new_n632), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n480), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n609), .A2(new_n242), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n620), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n407), .A2(new_n188), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n532), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT102), .Z(new_n644));
  NOR2_X1   g458(.A1(new_n475), .A2(KEYINPUT103), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n478), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n474), .A2(KEYINPUT103), .A3(new_n475), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n302), .A2(new_n650), .A3(new_n303), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n296), .A2(new_n300), .A3(KEYINPUT33), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n296), .A2(new_n300), .A3(KEYINPUT104), .A4(KEYINPUT33), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n305), .A2(G902), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n651), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n304), .A2(new_n305), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n262), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n644), .A2(new_n268), .A3(new_n649), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND2_X1  g478(.A1(new_n253), .A2(KEYINPUT20), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n251), .A2(new_n260), .A3(new_n252), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n304), .B(new_n310), .ZN(new_n668));
  INV_X1    g482(.A(new_n243), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n267), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n647), .A3(new_n646), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n644), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT105), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT35), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  INV_X1    g491(.A(new_n524), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n522), .A2(new_n481), .A3(new_n523), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n510), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n510), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n529), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT106), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n685), .A3(new_n529), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n679), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n527), .A2(KEYINPUT107), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n641), .A2(new_n642), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n316), .A2(new_n693), .A3(new_n479), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT37), .B(G110), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  NAND2_X1  g513(.A1(new_n624), .A2(new_n632), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n264), .B1(new_n265), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n670), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT107), .B1(new_n527), .B2(new_n688), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n524), .A2(new_n526), .A3(new_n690), .A4(new_n687), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n646), .A2(new_n188), .A3(new_n407), .A4(new_n647), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XNOR2_X1  g524(.A(new_n702), .B(KEYINPUT39), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n642), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT110), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n618), .A2(new_n606), .B1(new_n538), .B2(new_n586), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n614), .A2(new_n621), .A3(new_n622), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n476), .B(KEYINPUT38), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n262), .A2(new_n311), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n477), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n719), .A2(new_n693), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n714), .A2(new_n715), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  NOR3_X1   g538(.A1(new_n262), .A2(new_n660), .A3(new_n702), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n704), .B2(new_n705), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n707), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n700), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  AOI22_X1  g543(.A1(new_n373), .A2(new_n397), .B1(new_n401), .B2(new_n393), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n730), .B2(G902), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n405), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n188), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n527), .A3(new_n530), .ZN(new_n735));
  INV_X1    g549(.A(new_n262), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n659), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n648), .A2(new_n735), .A3(new_n737), .A4(new_n267), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n700), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  INV_X1    g555(.A(new_n735), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n700), .A2(new_n673), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  AND2_X1   g558(.A1(new_n316), .A2(new_n693), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n646), .A2(new_n647), .A3(new_n734), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n700), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n587), .A2(new_n537), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n619), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n605), .B(KEYINPUT111), .C1(new_n537), .C2(new_n587), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n608), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT112), .B(G472), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n753), .A2(new_n615), .B1(new_n639), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n531), .A2(new_n268), .A3(new_n755), .A4(new_n734), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n646), .A2(new_n720), .A3(new_n647), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(G122), .Z(G24));
  OAI21_X1  g573(.A(new_n755), .B1(new_n704), .B2(new_n705), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n725), .A2(new_n647), .A3(new_n646), .A4(new_n734), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n208), .ZN(G27));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n407), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n399), .A2(KEYINPUT113), .A3(new_n405), .A4(new_n406), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n188), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n476), .A2(new_n477), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n737), .A4(new_n702), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n629), .A2(new_n612), .A3(new_n621), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(KEYINPUT42), .A3(new_n531), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n633), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n772), .B1(new_n633), .B2(new_n769), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n771), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  NOR4_X1   g592(.A1(new_n767), .A2(new_n768), .A3(new_n670), .A4(new_n702), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n700), .A2(new_n779), .A3(new_n531), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  OR2_X1    g595(.A1(new_n398), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n398), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n406), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n406), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n785), .B(new_n405), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n188), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(new_n711), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT43), .B1(new_n262), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n262), .A2(new_n659), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n641), .A3(new_n693), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n768), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n792), .B(new_n799), .C1(new_n798), .C2(new_n797), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  XNOR2_X1  g615(.A(new_n790), .B(KEYINPUT47), .ZN(new_n802));
  INV_X1    g616(.A(new_n768), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n532), .A3(new_n725), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n700), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NOR3_X1   g620(.A1(new_n795), .A2(new_n733), .A3(new_n478), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n732), .A2(KEYINPUT49), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n531), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT117), .Z(new_n810));
  OAI21_X1  g624(.A(new_n719), .B1(KEYINPUT49), .B2(new_n732), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n810), .A2(new_n718), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n758), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n739), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n673), .A2(new_n742), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n316), .A2(new_n693), .A3(new_n746), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n816), .B1(new_n632), .B2(new_n624), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n667), .A2(new_n669), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n668), .A2(new_n702), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n768), .A2(new_n642), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n623), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n821), .B(new_n693), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n760), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n769), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n780), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n262), .A2(new_n659), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n311), .B2(new_n262), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n643), .A2(new_n829), .A3(new_n268), .A4(new_n479), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n695), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n637), .A2(new_n818), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n762), .B1(new_n700), .B2(new_n708), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n524), .A2(new_n526), .A3(new_n687), .A4(new_n702), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n718), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n757), .A3(new_n767), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n700), .B2(new_n727), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n834), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n838), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n833), .A2(new_n777), .A3(new_n842), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n846), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n833), .A2(new_n852), .A3(new_n853), .A4(new_n777), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n637), .A3(new_n832), .A4(new_n846), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n758), .B1(new_n700), .B2(new_n738), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n743), .A3(new_n747), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n747), .A3(new_n743), .A4(KEYINPUT120), .ZN(new_n861));
  AND4_X1   g675(.A1(KEYINPUT53), .A2(new_n780), .A3(new_n824), .A4(new_n826), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT54), .B1(new_n864), .B2(new_n777), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n842), .A2(new_n847), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n700), .A2(new_n531), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n635), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n633), .A2(KEYINPUT82), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n831), .B1(new_n870), .B2(new_n480), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n780), .A2(new_n824), .A3(new_n826), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n777), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n853), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n855), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n796), .A2(new_n264), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n531), .A3(new_n755), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n478), .A3(new_n719), .A4(new_n734), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT50), .Z(new_n881));
  OAI21_X1  g695(.A(new_n802), .B1(new_n188), .B2(new_n732), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n803), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n803), .A2(new_n734), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n531), .A2(new_n264), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n718), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n262), .A3(new_n660), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT121), .Z(new_n888));
  INV_X1    g702(.A(new_n884), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n878), .A2(new_n825), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(new_n883), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n878), .A2(new_n889), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n770), .A2(new_n531), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT48), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT122), .B(KEYINPUT48), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n879), .A2(new_n746), .ZN(new_n902));
  INV_X1    g716(.A(G952), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n903), .B(G953), .C1(new_n886), .C2(new_n661), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n899), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n877), .A2(new_n893), .A3(new_n894), .A4(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT123), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n812), .B1(new_n906), .B2(new_n908), .ZN(G75));
  AND3_X1   g723(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n777), .A3(new_n871), .A4(new_n852), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n875), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n444), .A2(new_n452), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n449), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT55), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n903), .A2(G953), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT124), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(G51));
  XOR2_X1   g737(.A(new_n406), .B(KEYINPUT57), .Z(new_n924));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n875), .A2(new_n925), .A3(new_n926), .A4(new_n911), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n848), .A2(new_n853), .B1(new_n864), .B2(new_n777), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n865), .B2(new_n875), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT126), .B(new_n924), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n403), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n912), .A2(G902), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(new_n784), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n922), .B1(new_n935), .B2(new_n937), .ZN(G54));
  NAND2_X1  g752(.A1(KEYINPUT58), .A2(G475), .ZN(new_n939));
  OR3_X1    g753(.A1(new_n936), .A2(new_n251), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n251), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n922), .B1(new_n940), .B2(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n855), .B2(new_n876), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n651), .A2(new_n655), .A3(new_n654), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n944), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n946), .B(new_n948), .C1(new_n929), .C2(new_n930), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n947), .A2(new_n921), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n928), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(new_n528), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n681), .A3(new_n682), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n921), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n921), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  NOR2_X1   g775(.A1(new_n447), .A2(new_n266), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n192), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n871), .A2(new_n818), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n192), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n915), .B1(G898), .B2(new_n192), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n965), .B(new_n966), .Z(G69));
  AND2_X1   g781(.A1(new_n834), .A2(new_n728), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n723), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT62), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n829), .A2(new_n803), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n713), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n870), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n805), .A2(new_n800), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n192), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n577), .A2(new_n578), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(new_n245), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n791), .A2(new_n757), .A3(new_n896), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n968), .A2(new_n780), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n974), .A2(new_n777), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n192), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n701), .A2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT127), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n979), .B1(new_n978), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n975), .B2(new_n964), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n537), .A3(new_n580), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n983), .B2(new_n964), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(new_n538), .A3(new_n576), .A4(new_n579), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n572), .B1(new_n601), .B2(new_n604), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n849), .A2(new_n854), .A3(new_n992), .A4(new_n997), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n921), .A2(new_n994), .A3(new_n996), .A4(new_n998), .ZN(G57));
endmodule


